VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO array_core
  CLASS BLOCK ;
  FOREIGN array_core ;
  ORIGIN 205.000 26.000 ;
  SIZE 609.600 BY 482.000 ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 127.000 443.000 135.000 456.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.000 443.000 49.000 456.000 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 61.000 448.000 69.000 456.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.000 -26.000 261.000 -24.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.000 448.000 155.000 456.000 ;
    END
  END VGND
  PIN a[0]
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 73.000 434.000 75.000 456.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 79.000 437.000 81.000 456.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 85.000 440.000 87.000 456.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 91.000 443.000 93.000 456.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 97.000 446.000 99.000 456.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 103.000 444.200 105.000 456.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 109.000 441.200 111.000 456.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 115.000 438.200 117.000 456.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.415000 ;
    PORT
      LAYER met3 ;
        RECT 121.000 435.200 123.000 456.000 ;
    END
  END a[8]
  PIN VTUN
    ANTENNADIFFAREA 759.539978 ;
    PORT
      LAYER met5 ;
        RECT 344.000 -26.000 366.000 -6.000 ;
    END
  END VTUN
  PIN VINJ
    ANTENNADIFFAREA 4575.179688 ;
    PORT
      LAYER met4 ;
        RECT 90.000 -26.000 110.000 -17.000 ;
    END
  END VINJ
  PIN VOUT0
    ANTENNADIFFAREA 15.080000 ;
    PORT
      LAYER met3 ;
        RECT 44.000 -26.000 48.000 -21.900 ;
    END
  END VOUT0
  PIN VCTRL
    ANTENNADIFFAREA 568.979980 ;
    PORT
      LAYER met3 ;
        RECT 28.600 -26.000 35.200 7.150 ;
    END
  END VCTRL
  PIN VSRC
    ANTENNADIFFAREA 174.000000 ;
    PORT
      LAYER met3 ;
        RECT 20.900 -26.000 27.500 -3.800 ;
    END
  END VSRC
  OBS
      LAYER nwell ;
        RECT -200.000 -18.000 399.830 446.230 ;
      LAYER li1 ;
        RECT -199.980 -17.670 399.810 446.210 ;
      LAYER met1 ;
        RECT -199.990 -22.000 399.820 446.220 ;
      LAYER met2 ;
        RECT -200.000 -22.000 402.420 446.230 ;
      LAYER met3 ;
        RECT -199.420 442.600 40.600 450.000 ;
        RECT 49.400 447.600 60.600 450.000 ;
        RECT 69.400 447.600 72.600 450.000 ;
        RECT 49.400 442.600 72.600 447.600 ;
        RECT -199.420 433.600 72.600 442.600 ;
        RECT 75.400 436.600 78.600 450.000 ;
        RECT 81.400 439.600 84.600 450.000 ;
        RECT 87.400 442.600 90.600 450.000 ;
        RECT 93.400 445.600 96.600 450.000 ;
        RECT 99.400 445.600 102.600 450.000 ;
        RECT 93.400 443.800 102.600 445.600 ;
        RECT 105.400 443.800 108.600 450.000 ;
        RECT 93.400 442.600 108.600 443.800 ;
        RECT 87.400 440.800 108.600 442.600 ;
        RECT 111.400 440.800 114.600 450.000 ;
        RECT 87.400 439.600 114.600 440.800 ;
        RECT 81.400 437.800 114.600 439.600 ;
        RECT 117.400 437.800 120.600 450.000 ;
        RECT 81.400 436.600 120.600 437.800 ;
        RECT 75.400 434.800 120.600 436.600 ;
        RECT 123.400 442.600 126.600 450.000 ;
        RECT 135.400 447.600 146.600 450.000 ;
        RECT 155.400 447.600 402.420 450.000 ;
        RECT 135.400 442.600 402.420 447.600 ;
        RECT 123.400 434.800 402.420 442.600 ;
        RECT 75.400 433.600 402.420 434.800 ;
        RECT -199.420 7.550 402.420 433.600 ;
        RECT -199.420 -3.400 28.200 7.550 ;
        RECT -199.420 -26.000 20.500 -3.400 ;
        RECT 27.900 -26.000 28.200 -3.400 ;
        RECT 35.600 -21.500 402.420 7.550 ;
        RECT 35.600 -26.000 43.600 -21.500 ;
        RECT 48.400 -23.600 402.420 -21.500 ;
        RECT 48.400 -26.000 238.600 -23.600 ;
        RECT 261.400 -26.000 402.420 -23.600 ;
      LAYER met4 ;
        RECT -205.000 -16.600 404.600 448.130 ;
        RECT -205.000 -23.000 89.600 -16.600 ;
        RECT 110.400 -23.000 404.600 -16.600 ;
      LAYER met5 ;
        RECT -205.000 -4.400 404.600 456.000 ;
        RECT -205.000 -15.000 342.400 -4.400 ;
        RECT 367.600 -15.000 404.600 -4.400 ;
  END
END array_core
END LIBRARY

