magic
tech sky130A
magscale 1 2
timestamp 1717473404
<< poly >>
rect 2907 -5477 3240 -5380
rect 3140 -5864 3240 -5477
rect 1336 -5964 3240 -5864
rect 3140 -6470 3240 -5964
<< locali >>
rect 3076 -5190 3282 -5060
<< metal1 >>
rect 3076 -5190 3322 -5098
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3360 -5194 3460 -5188
rect 4006 -7030 4106 -5098
rect 2900 -7130 4106 -7030
<< via1 >>
rect 3366 -5188 3454 -5100
rect 3508 -6552 3596 -6464
<< metal2 >>
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3360 -5222 3460 -5188
rect 2566 -5322 3460 -5222
rect 3502 -6464 3602 -6458
rect 3502 -6552 3508 -6464
rect 3596 -6552 3602 -6464
rect 3140 -6806 3240 -6770
rect 3502 -6806 3602 -6552
rect 1294 -6906 3602 -6806
use tg5v0  tg5v0_0
timestamp 1717473404
transform 0 -1 4094 1 0 -6628
box 28 0 1634 890
use fgcell  x1
timestamp 1717473404
transform 1 0 2010 0 1 -5490
box -1870 -310 1194 526
use diffamp_nmos  x2
timestamp 1717473404
transform 0 -1 3100 -1 0 -6070
box 20 -140 1140 2900
<< end >>
