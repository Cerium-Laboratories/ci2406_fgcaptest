magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< error_s >>
rect 2122 -5050 2442 -4980
rect 506 -5294 746 -5270
rect 506 -5486 530 -5294
rect 722 -5486 746 -5294
rect 2122 -5290 2146 -5050
rect 2372 -5290 2386 -5050
rect 2396 -5290 2442 -5050
rect 2122 -5314 2442 -5290
rect 506 -5510 746 -5486
rect 2992 -5501 3136 -5496
rect 2992 -5571 2997 -5501
rect 3131 -5571 3136 -5501
rect 2992 -5576 3136 -5571
rect 2506 -5651 2686 -5650
rect 2506 -5829 2507 -5651
rect 2685 -5829 2686 -5651
rect 2506 -5830 2686 -5829
rect 506 -6171 686 -6170
rect 506 -6349 507 -6171
rect 685 -6349 686 -6171
rect 3874 -6226 3880 -6220
rect 3920 -6226 3926 -6220
rect 3868 -6232 3874 -6226
rect 3926 -6232 3932 -6226
rect 3868 -6282 3874 -6276
rect 3926 -6282 3932 -6276
rect 3874 -6288 3880 -6282
rect 3920 -6288 3926 -6282
rect 506 -6350 686 -6349
rect 3402 -6402 3408 -6396
rect 3448 -6402 3454 -6396
rect 3396 -6408 3402 -6402
rect 3454 -6408 3460 -6402
rect 3396 -6454 3402 -6448
rect 3454 -6454 3460 -6448
rect 3402 -6460 3408 -6454
rect 3448 -6460 3454 -6454
rect 2526 -6914 2766 -6890
rect 2526 -7106 2550 -6914
rect 2742 -7106 2766 -6914
rect 2526 -7130 2766 -7106
<< poly >>
rect 2907 -5477 3240 -5380
rect 3140 -6470 3240 -5477
<< locali >>
rect 3076 -5190 3282 -5060
<< metal1 >>
rect 2136 -5050 2396 -5040
rect 2136 -5290 2146 -5050
rect 2386 -5290 2396 -5050
rect 2496 -5050 2656 -5040
rect 2496 -5190 2506 -5050
rect 2646 -5190 2656 -5050
rect 3076 -5190 3322 -5098
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 2496 -5200 2656 -5190
rect 3360 -5194 3460 -5188
rect 2136 -5300 2396 -5290
rect 3874 -6226 3932 -6220
rect 3926 -6282 3932 -6226
rect 3874 -6288 3932 -6282
rect 3396 -6402 3454 -6396
rect 3396 -6454 3402 -6402
rect 3396 -6458 3454 -6454
rect 3140 -6806 3240 -6670
rect 3502 -6806 3602 -6558
rect 3140 -6812 3602 -6806
rect 3234 -6900 3602 -6812
rect 3140 -6906 3602 -6900
rect 4006 -7030 4106 -5098
rect 2900 -7130 4106 -7030
<< via1 >>
rect 2146 -5290 2386 -5050
rect 2506 -5190 2646 -5050
rect 3366 -5188 3454 -5100
rect 3742 -5130 3830 -5042
rect 3874 -6282 3926 -6226
rect 3402 -6454 3454 -6402
rect 3140 -6900 3234 -6812
rect 410 -7104 896 -7036
rect 2586 -7130 2766 -7050
<< metal2 >>
rect 2136 -5050 2396 -5040
rect 496 -5270 756 -5260
rect 496 -5510 506 -5270
rect 746 -5510 756 -5270
rect 2136 -5290 2146 -5050
rect 2386 -5290 2396 -5050
rect 2496 -5050 2656 -5040
rect 2496 -5190 2506 -5050
rect 2646 -5190 2656 -5050
rect 3732 -5042 3840 -5032
rect 2496 -5200 2656 -5190
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3732 -5130 3742 -5042
rect 3830 -5130 3840 -5042
rect 3732 -5140 3840 -5130
rect 3360 -5222 3460 -5188
rect 2136 -5300 2396 -5290
rect 2706 -5322 3460 -5222
rect 496 -5520 756 -5510
rect 2758 -5496 3142 -5486
rect 2758 -5576 2992 -5496
rect 3136 -5576 3142 -5496
rect 2758 -5586 3142 -5576
rect 1294 -6812 3240 -6806
rect 1294 -6900 3140 -6812
rect 3234 -6900 3240 -6812
rect 496 -6910 696 -6900
rect 1294 -6906 3240 -6900
rect 496 -7030 506 -6910
rect 400 -7036 506 -7030
rect 686 -7030 696 -6910
rect 2576 -6950 2776 -6944
rect 686 -7036 906 -7030
rect 400 -7104 410 -7036
rect 896 -7104 906 -7036
rect 400 -7110 906 -7104
rect 2576 -7130 2586 -6950
rect 2766 -7130 2776 -6950
rect 2576 -7136 2776 -7130
<< via2 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2506 -5190 2646 -5050
rect 3742 -5130 3830 -5042
rect 2992 -5576 3136 -5496
rect 506 -7036 686 -6910
rect 506 -7090 686 -7036
rect 2586 -7050 2766 -6950
rect 2586 -7130 2766 -7050
<< metal3 >>
rect 2136 -5050 2396 -5040
rect 496 -5270 756 -5260
rect 496 -5510 506 -5270
rect 746 -5510 756 -5270
rect 2136 -5290 2146 -5050
rect 2386 -5290 2396 -5050
rect 2136 -5300 2396 -5290
rect 2486 -5050 2706 -5030
rect 2486 -5190 2506 -5050
rect 2646 -5190 2706 -5050
rect 3732 -5042 3840 -5032
rect 3732 -5130 3742 -5042
rect 3830 -5130 3840 -5042
rect 3732 -5140 3840 -5130
rect 496 -5520 756 -5510
rect 2486 -5650 2706 -5190
rect 2486 -5830 2506 -5650
rect 2686 -5830 2706 -5650
rect 2486 -5850 2706 -5830
rect 496 -6170 696 -6160
rect 496 -6350 506 -6170
rect 686 -6350 696 -6170
rect 496 -6910 696 -6350
rect 496 -7090 506 -6910
rect 686 -7090 696 -6910
rect 496 -7096 696 -7090
rect 2520 -6890 2776 -6884
rect 2520 -7130 2526 -6890
rect 2766 -7130 2776 -6890
rect 2520 -7140 2776 -7130
<< via3 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2506 -5830 2686 -5650
rect 506 -6350 686 -6170
rect 2526 -6950 2766 -6890
rect 2526 -7130 2586 -6950
rect 2586 -7130 2766 -6950
<< metal4 >>
rect 2136 -5050 2396 -5040
rect 496 -5270 756 -5260
rect 496 -5510 506 -5270
rect 746 -5510 756 -5270
rect 2136 -5290 2146 -5050
rect 2386 -5290 2396 -5050
rect 2136 -5300 2396 -5290
rect 496 -5520 756 -5510
rect 2520 -6890 2776 -6884
rect 2520 -7130 2526 -6890
rect 2766 -7130 2776 -6890
rect 2520 -7140 2776 -7130
<< via4 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2526 -7130 2766 -6890
<< metal5 >>
rect 2122 -5050 2396 -4980
rect 2122 -5290 2146 -5050
rect 2386 -5290 2396 -5050
rect 2122 -5314 2396 -5290
use tg5v0  tg5v0_0
timestamp 1717628967
transform 0 -1 4094 1 0 -6628
box 28 0 1634 890
use fgcell  x1
timestamp 1717628967
transform 1 0 2010 0 1 -5490
box -1870 -310 1194 526
use diffamp_nmos  x2
timestamp 1717628967
transform 0 -1 3100 -1 0 -6070
box 20 -140 1140 2900
<< labels >>
flabel metal3 3732 -5140 3840 -5032 0 FreeSans 32 0 0 0 vout
flabel metal1 3402 -6458 3454 -6402 0 FreeSans 160 0 0 0 row_en_b
flabel via1 3874 -6282 3926 -6226 0 FreeSans 160 0 0 0 row_en
flabel via4 2146 -5290 2386 -5050 0 FreeSans 320 0 0 0 VGND
flabel via4 2526 -7130 2766 -6890 0 FreeSans 640 0 0 0 VGND
flabel via2 2992 -5576 3136 -5496 0 FreeSans 320 0 0 0 VSRC
flabel via3 2506 -5830 2686 -5650 0 FreeSans 160 0 0 0 vinj
flabel via3 506 -6350 686 -6170 0 FreeSans 640 0 0 0 vdd
<< end >>
