magic
tech sky130A
magscale 1 2
timestamp 1717597221
<< nwell >>
rect -1704 198 -1174 322
rect -1704 28 -1136 198
rect -1704 -106 -1174 28
rect -670 -200 -84 416
rect 400 -248 1194 526
<< pwell >>
rect -1870 406 -1690 526
<< mvpmos >>
rect 697 168 897 268
rect -497 58 -297 158
rect 697 10 897 110
<< mvvaractor >>
rect -1487 58 -1287 158
<< mvpdiff >>
rect 697 314 897 326
rect 697 280 709 314
rect 885 280 897 314
rect 697 268 897 280
rect -497 204 -297 216
rect -497 170 -485 204
rect -309 170 -297 204
rect -497 158 -297 170
rect 697 110 897 168
rect -497 46 -297 58
rect -497 12 -485 46
rect -309 12 -297 46
rect -497 0 -297 12
rect 697 -2 897 10
rect 697 -36 709 -2
rect 885 -36 897 -2
rect 697 -48 897 -36
<< mvpdiffc >>
rect 709 280 885 314
rect -485 170 -309 204
rect -485 12 -309 46
rect 709 -36 885 -2
<< mvpsubdiff >>
rect -1870 506 -960 526
rect -1870 466 -1790 506
rect -1040 466 -960 506
rect -1870 446 -960 466
rect -1870 -230 -1790 446
rect -1040 392 -960 446
rect -1040 252 -1020 392
rect -980 252 -960 392
rect 160 392 240 416
rect -1040 228 -960 252
rect 160 252 180 392
rect 220 252 240 392
rect 160 228 240 252
rect -1040 -36 -960 -12
rect -1040 -176 -1020 -36
rect -980 -176 -960 -36
rect 160 -36 240 -12
rect -1040 -230 -960 -176
rect 160 -176 180 -36
rect 220 -176 240 -36
rect 160 -200 240 -176
rect -1870 -250 -960 -230
rect -1870 -290 -1790 -250
rect -1040 -290 -960 -250
rect -1870 -310 -960 -290
<< mvnsubdiff >>
rect 466 448 1066 460
rect -1487 243 -1287 255
rect -1487 220 -1463 243
rect -1638 209 -1463 220
rect -1311 209 -1287 243
rect 466 414 574 448
rect 1020 414 1066 448
rect 466 402 1066 414
rect -604 338 -150 350
rect -604 304 -580 338
rect -174 304 -150 338
rect -604 292 -150 304
rect -1638 196 -1287 209
rect -1638 82 -1632 196
rect -1598 176 -1287 196
rect -1598 82 -1594 176
rect -1487 158 -1287 176
rect -1638 58 -1594 82
rect -1487 7 -1287 58
rect -1487 -27 -1463 7
rect -1311 -27 -1287 7
rect -1487 -39 -1287 -27
rect -604 -88 -150 -76
rect -604 -122 -580 -88
rect -174 -122 -150 -88
rect -604 -134 -150 -122
rect 466 -136 1066 -124
rect 466 -170 574 -136
rect 1020 -170 1066 -136
rect 466 -182 1066 -170
<< mvpsubdiffcont >>
rect -1790 466 -1040 506
rect -1020 252 -980 392
rect 180 252 220 392
rect -1020 -176 -980 -36
rect 180 -176 220 -36
rect -1790 -290 -1040 -250
<< mvnsubdiffcont >>
rect -1463 209 -1311 243
rect 574 414 1020 448
rect -580 304 -174 338
rect -1632 82 -1598 196
rect -1463 -27 -1311 7
rect -580 -122 -174 -88
rect 574 -170 1020 -136
<< poly >>
rect 656 168 697 268
rect 897 252 994 268
rect 897 184 944 252
rect 978 184 994 252
rect 897 168 994 184
rect -1575 58 -1487 158
rect -1287 142 -1166 158
rect -1287 74 -1248 142
rect -1176 74 -1166 142
rect -1287 58 -1166 74
rect -1124 142 -497 158
rect -1124 74 -1114 142
rect -1042 74 -497 142
rect -1124 58 -497 74
rect -297 110 500 158
rect -297 58 697 110
rect 400 10 697 58
rect 897 10 994 110
<< polycont >>
rect 944 184 978 252
rect -1248 74 -1176 142
rect -1114 74 -1042 142
<< locali >>
rect -1866 512 -964 522
rect -1866 454 -1856 512
rect -1798 506 -964 512
rect -1798 466 -1790 506
rect -1040 466 -964 506
rect -1798 454 -964 466
rect -1866 450 -964 454
rect -1866 392 -1794 450
rect -1866 -176 -1850 392
rect -1810 -176 -1794 392
rect -1036 392 -964 450
rect 478 414 574 448
rect 1020 414 1066 448
rect -1036 252 -1020 392
rect -980 252 -964 392
rect -604 304 -580 338
rect -174 304 -150 338
rect 164 252 180 392
rect 220 252 236 392
rect 478 314 1066 414
rect 478 302 709 314
rect 693 280 709 302
rect 885 302 1066 314
rect 885 280 901 302
rect 944 252 978 268
rect -1632 243 -1294 244
rect -1632 209 -1463 243
rect -1311 209 -1294 243
rect -1632 208 -1294 209
rect -1632 196 -1598 208
rect -501 170 -485 204
rect -309 170 -293 204
rect 944 168 978 184
rect -1632 66 -1598 82
rect -1264 74 -1248 142
rect -1176 74 -1114 142
rect -1042 74 -1026 142
rect -501 12 -485 46
rect -309 12 -293 46
rect -1479 -27 -1463 7
rect -1311 -27 -1295 7
rect 693 -36 709 -2
rect 885 -36 901 -2
rect -1866 -234 -1794 -176
rect -1036 -176 -1020 -36
rect -980 -176 -964 -36
rect -604 -122 -580 -88
rect -174 -122 -150 -88
rect 164 -176 180 -36
rect 220 -176 236 -36
rect 478 -170 574 -136
rect 1020 -170 1066 -136
rect -1036 -234 -964 -176
rect -1866 -250 -964 -234
rect -1866 -290 -1790 -250
rect -1040 -290 -964 -250
rect -1866 -306 -964 -290
<< viali >>
rect -1856 454 -1798 512
rect -1700 466 -1040 506
rect -1850 -176 -1810 392
rect 574 414 1020 448
rect -1020 252 -980 392
rect -580 304 -174 338
rect 180 252 220 392
rect 709 280 885 314
rect -1463 209 -1311 243
rect -1632 82 -1598 196
rect -485 170 -309 204
rect 944 184 978 252
rect -485 12 -309 46
rect -1463 -27 -1311 7
rect 709 -36 885 -2
rect -1020 -176 -980 -36
rect -580 -122 -174 -88
rect 180 -176 220 -36
rect 574 -170 1020 -136
rect -1790 -290 -1040 -250
<< metal1 >>
rect -1868 518 236 524
rect -1868 434 -1862 518
rect -1778 506 236 518
rect -1778 466 -1700 506
rect -1040 466 236 506
rect -1778 450 236 466
rect -1778 434 -1772 450
rect -1868 428 -1772 434
rect -1868 392 -1794 428
rect -1868 -176 -1850 392
rect -1810 -176 -1794 392
rect -1036 392 -964 450
rect -1036 252 -1020 392
rect -980 252 -964 392
rect 164 392 236 450
rect -592 338 -162 344
rect -592 304 -580 338
rect -174 304 -162 338
rect -592 298 -162 304
rect -1638 244 -1298 250
rect -1036 246 -964 252
rect -1638 243 -1456 244
rect -1318 243 -1298 244
rect -1638 209 -1463 243
rect -1311 209 -1298 243
rect -452 210 -352 298
rect 164 252 180 392
rect 220 252 236 392
rect -1638 202 -1456 209
rect -1638 196 -1592 202
rect -1638 82 -1632 196
rect -1598 82 -1592 196
rect -1638 70 -1592 82
rect -1463 192 -1456 202
rect -1318 202 -1298 209
rect -497 204 -297 210
rect -1318 192 -1311 202
rect -1463 24 -1311 192
rect -497 170 -485 204
rect -309 170 -297 204
rect -497 164 -297 170
rect -452 52 -352 164
rect -1463 13 -1456 24
rect -1475 7 -1456 13
rect -1318 13 -1311 24
rect -497 46 -297 52
rect -1318 7 -1299 13
rect -1475 -27 -1463 7
rect -1311 -27 -1299 7
rect -497 12 -485 46
rect -309 12 -297 46
rect -497 6 -297 12
rect -1475 -28 -1456 -27
rect -1318 -28 -1299 -27
rect -1475 -33 -1299 -28
rect -1868 -234 -1794 -176
rect -1036 -36 -964 -30
rect -1036 -176 -1020 -36
rect -980 -176 -964 -36
rect -452 -82 -352 6
rect 164 -36 236 252
rect -592 -88 -162 -82
rect -592 -122 -580 -88
rect -174 -122 -162 -88
rect -592 -128 -162 -122
rect -1036 -234 -964 -176
rect -1868 -250 -964 -234
rect -1868 -290 -1790 -250
rect -1040 -290 -964 -250
rect -1868 -306 -964 -290
rect -452 -204 -352 -128
rect 164 -176 180 -36
rect 220 -176 236 -36
rect 478 448 1066 454
rect 478 414 574 448
rect 1020 414 1066 448
rect 478 396 1066 414
rect 478 336 806 396
rect 478 -130 638 336
rect 696 314 806 336
rect 890 336 1066 396
rect 696 280 709 314
rect 890 312 898 336
rect 885 280 898 312
rect 696 274 898 280
rect 938 260 1038 268
rect 938 252 946 260
rect 938 184 944 252
rect 938 176 946 184
rect 1030 176 1038 260
rect 938 168 1038 176
rect 697 -2 897 4
rect 697 -36 709 -2
rect 885 -36 897 -2
rect 697 -42 756 -36
rect 748 -88 756 -42
rect 840 -42 897 -36
rect 840 -88 848 -42
rect 748 -96 848 -88
rect 478 -136 1066 -130
rect 478 -170 574 -136
rect 1020 -170 1066 -136
rect 478 -176 1066 -170
rect 164 -182 236 -176
rect -452 -288 -444 -204
rect -360 -288 -352 -204
rect -452 -296 -352 -288
<< via1 >>
rect -1862 512 -1778 518
rect -1862 454 -1856 512
rect -1856 454 -1798 512
rect -1798 454 -1778 512
rect -1862 434 -1778 454
rect -1456 243 -1318 244
rect -1456 209 -1318 243
rect -1456 192 -1318 209
rect -1456 7 -1318 24
rect -1456 -27 -1318 7
rect -1456 -28 -1318 -27
rect 806 314 890 396
rect 806 312 885 314
rect 885 312 890 314
rect 946 252 1030 260
rect 946 184 978 252
rect 978 184 1030 252
rect 946 176 1030 184
rect 756 -36 840 -4
rect 756 -88 840 -36
rect -444 -288 -360 -204
<< metal2 >>
rect -1870 518 -1770 526
rect -1870 434 -1862 518
rect -1778 434 -1770 518
rect -1870 426 -1770 434
rect 798 396 898 404
rect 798 312 806 396
rect 890 312 898 396
rect 798 304 898 312
rect 938 260 1038 268
rect -1462 192 -1456 244
rect -1318 192 -1312 244
rect -1462 24 -1312 192
rect 938 176 946 260
rect 1030 176 1038 260
rect 938 168 1038 176
rect -1462 -28 -1456 24
rect -1318 -28 -1312 24
rect 748 -4 848 4
rect 748 -88 756 -4
rect 840 -88 848 -4
rect 748 -96 848 -88
rect -452 -204 -352 -196
rect -452 -288 -444 -204
rect -360 -288 -352 -204
rect -452 -296 -352 -288
<< labels >>
flabel poly -1104 58 -1054 158 0 FreeSans 480 0 0 0 fg
flabel metal2 -452 -296 -352 -196 0 FreeSans 480 0 0 0 vctrl
port 3 nsew analog input
flabel metal2 748 -96 848 4 0 FreeSans 480 0 0 0 vsrc
port 4 nsew signal input
flabel metal2 798 304 898 404 0 FreeSans 480 0 0 0 vinj
port 0 nsew power default
flabel poly -6 58 94 158 0 FreeSans 320 0 0 0 vfg
port 6 nsew
flabel metal2 -1870 426 -1770 526 0 FreeSans 480 0 0 0 VGND
port 5 nsew ground default
flabel metal2 -1462 -28 -1312 244 0 FreeSans 480 0 0 0 vtun
port 2 nsew analog input
flabel metal2 938 168 1038 268 0 FreeSans 480 180 0 0 vinj_en_b
port 1 nsew signal input
<< properties >>
string FIXED_BBOX -2010 -510 1394 726
<< end >>
