* NGSPICE file created from diffamp_nmos.ext - technology: sky130A

.subckt diffamp_nmos v1 v2 VSS VDD vb vout
X0 a_400_700# vb int1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X1 int3 int3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X2 VSS vb a_400_700# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X3 int1 v1 int4 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X4 VDD int4 int4 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X5 VSS int2 int2 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X6 int3 v2 int1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X7 vout int2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X8 VDD int3 int2 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X9 vout int4 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
.ends

