** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/test-fgcell.sch
**.subckt test-fgcell
x1 vinj vinj_en_b vfg vtun vctrl vsrc GND fgcell
vinj_en_b vinj_en_b GND pwl(0 {VINJ} 80u {VINJ} 85u 0)
vctrl vctrl GND 0 pwl(0 0 10u 0 15u {VINJ} 20u {VINJ} 25u 0)
vsrc vsrc GND pwl(0 {VINJ} 70u {VINJ} 75u 0)
vtun vtun GND pwl(0 0 30u 0 40u {VTUN} 50u {VTUN} 60u 0)
vinj vinj GND {VINJ}
R1 vfg GND 1T m=1
**** begin user architecture code
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.options reltol=0.0001 abstol=10e-15 chgtol=1e-15
* .include fgcell.spice
.param VTUN=12
.param VINJ=6
.param VDD=1.8
.param VSS=0
.option savecurrents
.ic v(vinj)=6 v(vinj_en_b)=6 v(vtun)=0 v(vsrc)=6 v(vfg)=0 v(x1.net1)=6
.control
  save all
  *op
  *remzerovec
  *write test-fgcell.raw
  *set appendwrite
  tran 10n 120u uic
  remzerovec
  write test-fgcell.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  fgcell.sym # of pins=7
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/fgcell.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/fgcell.sch
.subckt fgcell vinj vinj_en_b vfg vtun vctrl vsrc VGND
*.ipin vctrl
*.ipin vtun
*.ipin vinj
*.ipin vinj_en_b
*.ipin vsrc
*.opin vfg
*.ipin VGND
XC1 vfg vtun vtun sky130_fd_pr__cap_var_hvt W=0.5 L=0.5 VM=1 m=1
XM1 vsrc vfg net1 vinj sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 vinj_en_b vinj vinj sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vctrl vfg vctrl vctrl sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
