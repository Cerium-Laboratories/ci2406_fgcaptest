magic
tech sky130A
magscale 1 2
timestamp 1717346353
<< error_p >>
rect 37560 12304 37680 12310
rect 37588 12276 37652 12282
rect 9770 -13600 9783 -13364
rect 20219 -13380 20243 -13364
rect 20243 -13600 20246 -13380
rect 54770 -13600 54783 -13380
rect 80219 -13380 80243 -13364
rect 80243 -13600 80246 -13380
rect 9451 -13688 9684 -13672
rect 9448 -13908 9451 -13688
rect 20372 -13742 20605 -13726
rect 20605 -13962 20608 -13742
rect 65372 -13742 65551 -13726
rect 54448 -13908 54451 -13742
rect 80372 -13742 80605 -13726
rect 80605 -13962 80608 -13742
rect 9141 -13998 9364 -13992
rect 9128 -14228 9141 -13998
rect 20692 -14056 20919 -14046
rect 20919 -14282 20928 -14056
rect 65692 -14056 65861 -14046
rect 54128 -14228 54141 -14056
rect 80692 -14056 80919 -14046
rect 80919 -14282 80928 -14056
rect 8811 -14328 9044 -14312
rect 8808 -14548 8811 -14328
rect 21012 -14382 21240 -14366
rect 66012 -14382 66191 -14366
rect 53808 -14548 53811 -14382
rect 81012 -14382 81245 -14366
rect 81245 -14390 81248 -14382
rect 8497 -14642 8721 -14635
rect 8485 -14662 8497 -14642
rect 9943 -21517 9977 -21483
rect 9979 -21555 10015 -21483
rect 8754 -27378 8757 -27158
rect 8757 -27394 8990 -27378
rect 9074 -27698 9077 -27478
rect 9077 -27714 9310 -27698
rect 9394 -28018 9397 -27798
rect 9397 -28034 9630 -28018
rect 9756 -28380 9759 -28160
rect 9759 -28396 9783 -28380
<< error_s >>
rect 53356 -8776 53412 -8720
rect 24770 -13600 24783 -13364
rect 35219 -13380 35243 -13364
rect 35243 -13600 35246 -13380
rect 24451 -13688 24684 -13672
rect 24448 -13908 24451 -13688
rect 35551 -13742 35605 -13726
rect 35605 -13962 35608 -13742
rect 24141 -13998 24364 -13992
rect 24128 -14228 24141 -13998
rect 35861 -14056 35919 -14046
rect 35919 -14282 35928 -14056
rect 23811 -14328 24044 -14312
rect 21240 -14382 21245 -14366
rect 23808 -14373 23811 -14328
rect 36191 -14382 36245 -14366
rect 21245 -14390 21248 -14382
rect 36245 -14390 36248 -14382
rect 51240 -14382 51245 -14366
rect 66240 -14382 66245 -14366
rect 51245 -14390 51248 -14382
rect 66245 -14390 66248 -14382
rect 23497 -14642 23721 -14635
rect 38497 -14642 38721 -14635
rect 53497 -14642 53721 -14635
rect 68497 -14642 68721 -14635
rect 23485 -14662 23497 -14642
rect 38485 -14662 38497 -14642
rect 53485 -14662 53497 -14642
rect 68485 -14662 68497 -14642
rect 19985 -21555 20021 -21483
rect 20023 -21517 20057 -21483
rect 24943 -21517 24977 -21483
rect 24979 -21555 25015 -21483
rect 34985 -21555 35021 -21483
rect 35023 -21517 35057 -21483
rect 39943 -21517 39977 -21483
rect 39979 -21555 40015 -21483
rect 49985 -21555 50021 -21483
rect 50023 -21517 50057 -21483
rect 54943 -21517 54977 -21483
rect 54979 -21555 55015 -21483
rect 64985 -21555 65021 -21483
rect 65023 -21517 65057 -21483
rect 69943 -21517 69977 -21483
rect 69979 -21555 70015 -21483
rect 79985 -21555 80021 -21483
rect 80023 -21517 80057 -21483
rect 21514 -27109 21517 -27098
rect 36514 -27109 36517 -27098
rect 51514 -27109 51517 -27098
rect 66514 -27109 66517 -27098
rect 81514 -27109 81517 -27098
rect 21286 -27125 21514 -27109
rect 36286 -27125 36514 -27109
rect 51286 -27125 51514 -27109
rect 66286 -27125 66514 -27109
rect 81286 -27125 81514 -27109
rect 23754 -27378 23757 -27337
rect 38754 -27378 38757 -27158
rect 53754 -27378 53757 -27337
rect 68754 -27378 68757 -27158
rect 21191 -27432 21194 -27380
rect 23757 -27387 23766 -27378
rect 23766 -27394 23990 -27387
rect 36191 -27432 36194 -27380
rect 38757 -27394 38990 -27378
rect 53757 -27380 53759 -27378
rect 51191 -27432 51194 -27380
rect 53759 -27394 53811 -27380
rect 66191 -27432 66194 -27380
rect 68757 -27394 68990 -27378
rect 81191 -27432 81194 -27380
rect 20958 -27448 21191 -27432
rect 35958 -27448 36191 -27432
rect 50958 -27448 51191 -27432
rect 65958 -27448 66191 -27432
rect 80958 -27448 81191 -27432
rect 20871 -27752 20874 -27532
rect 24074 -27698 24077 -27478
rect 39074 -27698 39077 -27478
rect 24077 -27714 24310 -27698
rect 35871 -27752 35874 -27698
rect 39077 -27714 39310 -27698
rect 50871 -27752 50874 -27532
rect 54074 -27698 54077 -27478
rect 69074 -27698 69077 -27478
rect 54077 -27714 54131 -27698
rect 65871 -27752 65874 -27698
rect 69077 -27714 69310 -27698
rect 80871 -27752 80874 -27532
rect 20754 -27768 20871 -27752
rect 35754 -27768 35871 -27752
rect 50754 -27768 50871 -27752
rect 65754 -27768 65871 -27752
rect 80754 -27768 80871 -27752
rect 20551 -28072 20554 -27869
rect 24394 -28018 24397 -27798
rect 39394 -28018 39397 -27798
rect 24397 -28034 24630 -28018
rect 35551 -28072 35554 -28018
rect 39397 -28034 39630 -28018
rect 50551 -28072 50554 -27869
rect 54394 -28018 54397 -27869
rect 69394 -28018 69397 -27798
rect 54397 -28034 54451 -28018
rect 65551 -28072 65554 -28018
rect 69397 -28034 69630 -28018
rect 80551 -28072 80554 -27869
rect 20318 -28088 20551 -28072
rect 35318 -28088 35551 -28072
rect 50318 -28088 50551 -28072
rect 65318 -28088 65551 -28072
rect 80318 -28088 80551 -28072
rect 20219 -28396 20232 -28160
rect 24756 -28380 24759 -28160
rect 39756 -28380 39759 -28160
rect 24759 -28396 24783 -28380
rect 35219 -28396 35232 -28380
rect 39759 -28396 39783 -28380
rect 50219 -28396 50232 -28160
rect 54756 -28380 54759 -28160
rect 69756 -28380 69759 -28160
rect 54759 -28396 54783 -28380
rect 65219 -28396 65232 -28380
rect 69759 -28396 69783 -28380
rect 80219 -28396 80232 -28160
<< error_ps >>
rect 39770 -13600 39783 -13364
rect 50219 -13380 50243 -13364
rect 54770 -13380 54783 -13364
rect 65219 -13380 65243 -13364
rect 50243 -13600 50246 -13380
rect 65243 -13600 65246 -13380
rect 69770 -13600 69783 -13364
rect 39451 -13688 39684 -13672
rect 54451 -13688 54684 -13672
rect 69451 -13688 69684 -13672
rect 39448 -13908 39451 -13688
rect 50372 -13742 50605 -13726
rect 54448 -13742 54451 -13688
rect 65551 -13742 65605 -13726
rect 50605 -13962 50608 -13742
rect 65605 -13962 65608 -13742
rect 69448 -13908 69451 -13688
rect 39141 -13998 39364 -13992
rect 54141 -13998 54364 -13992
rect 69141 -13998 69364 -13992
rect 39128 -14228 39141 -13998
rect 50692 -14056 50919 -14046
rect 54128 -14056 54141 -13998
rect 65861 -14056 65919 -14046
rect 50919 -14282 50928 -14056
rect 65919 -14282 65928 -14056
rect 69128 -14228 69141 -13998
rect 38811 -14328 39044 -14312
rect 53811 -14328 54044 -14312
rect 68811 -14328 69044 -14312
rect 38808 -14548 38811 -14328
rect 51012 -14382 51240 -14366
rect 53808 -14382 53811 -14328
rect 66191 -14382 66240 -14366
rect 68808 -14548 68811 -14328
<< metal1 >>
rect 64882 3960 65038 3966
rect 51996 3954 64882 3960
rect 51996 3902 52028 3954
rect 52132 3902 53628 3954
rect 53732 3902 55228 3954
rect 55332 3902 56828 3954
rect 56932 3902 58428 3954
rect 58532 3902 60028 3954
rect 60132 3902 61628 3954
rect 61732 3902 63228 3954
rect 63332 3902 64882 3954
rect 51996 3800 64882 3902
rect 52360 3708 52476 3714
rect 52360 3604 52366 3708
rect 52470 3604 52476 3708
rect 52746 3688 52830 3800
rect 53160 3708 53276 3714
rect 52360 3598 52476 3604
rect 53160 3604 53166 3708
rect 53270 3604 53276 3708
rect 53546 3688 53630 3800
rect 53960 3708 54076 3714
rect 53160 3598 53276 3604
rect 53960 3604 53966 3708
rect 54070 3604 54076 3708
rect 54346 3688 54430 3800
rect 54760 3708 54876 3714
rect 53960 3598 54076 3604
rect 54760 3604 54766 3708
rect 54870 3604 54876 3708
rect 55146 3688 55230 3800
rect 55560 3708 55676 3714
rect 54760 3598 54876 3604
rect 55560 3604 55566 3708
rect 55670 3604 55676 3708
rect 55946 3688 56030 3800
rect 56360 3708 56476 3714
rect 55560 3598 55676 3604
rect 56360 3604 56366 3708
rect 56470 3604 56476 3708
rect 56746 3688 56830 3800
rect 57160 3708 57276 3714
rect 56360 3598 56476 3604
rect 57160 3604 57166 3708
rect 57270 3604 57276 3708
rect 57546 3688 57630 3800
rect 57960 3708 58076 3714
rect 57160 3598 57276 3604
rect 57960 3604 57966 3708
rect 58070 3604 58076 3708
rect 58346 3688 58430 3800
rect 58760 3708 58876 3714
rect 57960 3598 58076 3604
rect 58760 3604 58766 3708
rect 58870 3604 58876 3708
rect 59146 3688 59230 3800
rect 59560 3708 59676 3714
rect 58760 3598 58876 3604
rect 59560 3604 59566 3708
rect 59670 3604 59676 3708
rect 59946 3688 60030 3800
rect 60360 3708 60476 3714
rect 59560 3598 59676 3604
rect 60360 3604 60366 3708
rect 60470 3604 60476 3708
rect 60746 3688 60830 3800
rect 61160 3708 61276 3714
rect 60360 3598 60476 3604
rect 61160 3604 61166 3708
rect 61270 3604 61276 3708
rect 61546 3688 61630 3800
rect 61960 3708 62076 3714
rect 61160 3598 61276 3604
rect 61960 3604 61966 3708
rect 62070 3604 62076 3708
rect 62346 3688 62430 3800
rect 62760 3708 62876 3714
rect 61960 3598 62076 3604
rect 62760 3604 62766 3708
rect 62870 3604 62876 3708
rect 63146 3688 63230 3800
rect 63560 3708 63676 3714
rect 62760 3598 62876 3604
rect 63560 3604 63566 3708
rect 63670 3604 63676 3708
rect 63946 3688 64030 3800
rect 64360 3708 64476 3714
rect 63560 3598 63676 3604
rect 64360 3604 64366 3708
rect 64470 3604 64476 3708
rect 64746 3688 64830 3800
rect 64882 3794 65038 3800
rect 64360 3598 64476 3604
<< via1 >>
rect 52028 4260 52132 4312
rect 53628 4260 53732 4312
rect 55228 4260 55332 4312
rect 56828 4260 56932 4312
rect 58428 4260 58532 4312
rect 60028 4260 60132 4312
rect 61628 4260 61732 4312
rect 63228 4260 63332 4312
rect 52028 3902 52132 3954
rect 53628 3902 53732 3954
rect 55228 3902 55332 3954
rect 56828 3902 56932 3954
rect 58428 3902 58532 3954
rect 60028 3902 60132 3954
rect 61628 3902 61732 3954
rect 63228 3902 63332 3954
rect 64882 3800 65038 3960
rect 52366 3604 52470 3708
rect 53166 3604 53270 3708
rect 53966 3604 54070 3708
rect 54766 3604 54870 3708
rect 55566 3604 55670 3708
rect 56366 3604 56470 3708
rect 57166 3604 57270 3708
rect 57966 3604 58070 3708
rect 58766 3604 58870 3708
rect 59566 3604 59670 3708
rect 60366 3604 60470 3708
rect 61166 3604 61270 3708
rect 61966 3604 62070 3708
rect 62766 3604 62870 3708
rect 63566 3604 63670 3708
rect 64366 3604 64470 3708
<< metal2 >>
rect 52022 4312 52138 4318
rect 52022 4260 52028 4312
rect 52132 4260 52138 4312
rect 52022 3954 52138 4260
rect 53622 4312 53738 4318
rect 53622 4260 53628 4312
rect 53732 4260 53738 4312
rect 52022 3902 52028 3954
rect 52132 3902 52138 3954
rect 52022 3896 52138 3902
rect 52360 3708 52476 4000
rect 52360 3604 52366 3708
rect 52470 3604 52476 3708
rect 52360 3598 52476 3604
rect 53160 3708 53276 4000
rect 53622 3954 53738 4260
rect 55222 4312 55338 4318
rect 55222 4260 55228 4312
rect 55332 4260 55338 4312
rect 53622 3902 53628 3954
rect 53732 3902 53738 3954
rect 53622 3896 53738 3902
rect 53160 3604 53166 3708
rect 53270 3604 53276 3708
rect 53160 3598 53276 3604
rect 53960 3708 54076 4000
rect 53960 3604 53966 3708
rect 54070 3604 54076 3708
rect 53960 3598 54076 3604
rect 54760 3708 54876 4000
rect 55222 3954 55338 4260
rect 56822 4312 56938 4318
rect 56822 4260 56828 4312
rect 56932 4260 56938 4312
rect 55222 3902 55228 3954
rect 55332 3902 55338 3954
rect 55222 3896 55338 3902
rect 54760 3604 54766 3708
rect 54870 3604 54876 3708
rect 54760 3598 54876 3604
rect 55560 3708 55676 4000
rect 55560 3604 55566 3708
rect 55670 3604 55676 3708
rect 55560 3598 55676 3604
rect 56360 3708 56476 4000
rect 56822 3954 56938 4260
rect 58422 4312 58538 4318
rect 58422 4260 58428 4312
rect 58532 4260 58538 4312
rect 56822 3902 56828 3954
rect 56932 3902 56938 3954
rect 56822 3896 56938 3902
rect 56360 3604 56366 3708
rect 56470 3604 56476 3708
rect 56360 3598 56476 3604
rect 57160 3708 57276 4000
rect 57160 3604 57166 3708
rect 57270 3604 57276 3708
rect 57160 3598 57276 3604
rect 57960 3708 58076 4000
rect 58422 3954 58538 4260
rect 60022 4312 60138 4318
rect 60022 4260 60028 4312
rect 60132 4260 60138 4312
rect 58422 3902 58428 3954
rect 58532 3902 58538 3954
rect 58422 3896 58538 3902
rect 57960 3604 57966 3708
rect 58070 3604 58076 3708
rect 57960 3598 58076 3604
rect 58760 3708 58876 4000
rect 58760 3604 58766 3708
rect 58870 3604 58876 3708
rect 58760 3598 58876 3604
rect 59560 3708 59676 4000
rect 60022 3954 60138 4260
rect 61622 4312 61738 4318
rect 61622 4260 61628 4312
rect 61732 4260 61738 4312
rect 60022 3902 60028 3954
rect 60132 3902 60138 3954
rect 60022 3896 60138 3902
rect 59560 3604 59566 3708
rect 59670 3604 59676 3708
rect 59560 3598 59676 3604
rect 60360 3708 60476 4000
rect 60360 3604 60366 3708
rect 60470 3604 60476 3708
rect 60360 3598 60476 3604
rect 61160 3708 61276 4000
rect 61622 3954 61738 4260
rect 63222 4312 63338 4318
rect 63222 4260 63228 4312
rect 63332 4260 63338 4312
rect 61622 3902 61628 3954
rect 61732 3902 61738 3954
rect 61622 3896 61738 3902
rect 61160 3604 61166 3708
rect 61270 3604 61276 3708
rect 61160 3598 61276 3604
rect 61960 3708 62076 4000
rect 61960 3604 61966 3708
rect 62070 3604 62076 3708
rect 61960 3598 62076 3604
rect 62760 3708 62876 4000
rect 63222 3954 63338 4260
rect 63222 3902 63228 3954
rect 63332 3902 63338 3954
rect 63222 3896 63338 3902
rect 62760 3604 62766 3708
rect 62870 3604 62876 3708
rect 62760 3598 62876 3604
rect 63560 3708 63676 4000
rect 63560 3604 63566 3708
rect 63670 3604 63676 3708
rect 63560 3598 63676 3604
rect 64360 3708 64476 4000
rect 64882 3960 65038 4260
rect 64882 3794 65038 3800
rect 64360 3604 64366 3708
rect 64470 3604 64476 3708
rect 64360 3598 64476 3604
<< metal3 >>
rect 50200 89800 51800 90000
rect 52200 89800 53800 90000
rect 54600 89800 55000 90000
rect 55800 89800 56200 90000
rect 57000 89800 57400 90000
rect 58200 89800 58600 90000
rect 59400 89800 59800 90000
rect 60600 89800 61000 90000
rect 61800 89800 62200 90000
rect 63000 89800 63400 90000
rect 64200 89800 64600 90000
rect 65400 89800 67000 90000
rect 67400 89800 69000 90000
use array_core  array_core_0
timestamp 1717346353
transform 1 0 40000 0 1 0
box -40000 -3600 79966 90000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1717304525
transform -1 0 37500 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_1
timestamp 1717304525
transform -1 0 22500 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_2
timestamp 1717304525
transform -1 0 67500 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_3
timestamp 1717304525
transform -1 0 52500 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_4
timestamp 1717304525
transform -1 0 82500 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1717304525
transform 1 0 105000 0 1 -27880
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_2
timestamp 1717304525
transform 1 0 84000 0 1 -27880
box -540 -540 12540 14540
<< labels >>
flabel metal3 50200 89800 51800 90000 0 FreeSans 1600 0 0 0 vccd1
port 1 nsew power default
flabel metal3 52200 89800 53800 90000 0 FreeSans 1600 0 0 0 vssd1
port 2 nsew ground default
flabel metal3 54600 89800 55000 90000 0 FreeSans 800 0 0 0 addr[0]
port 3 nsew signal input
flabel metal3 55800 89800 56200 90000 0 FreeSans 800 0 0 0 addr[1]
port 4 nsew signal input
flabel metal3 57000 89800 57400 90000 0 FreeSans 800 0 0 0 addr[2]
port 5 nsew signal input
flabel metal3 58200 89800 58600 90000 0 FreeSans 800 0 0 0 addr[3]
port 6 nsew signal input
flabel metal3 59400 89800 59800 90000 0 FreeSans 800 0 0 0 addr[4]
port 7 nsew signal input
flabel metal3 60600 89800 61000 90000 0 FreeSans 800 0 0 0 addr[5]
port 8 nsew signal input
flabel metal3 61800 89800 62200 90000 0 FreeSans 800 0 0 0 addr[6]
port 9 nsew signal input
flabel metal3 63000 89800 63400 90000 0 FreeSans 800 0 0 0 addr[7]
port 10 nsew signal input
flabel metal3 64200 89800 64600 90000 0 FreeSans 800 0 0 0 addr[8]
port 11 nsew signal input
flabel metal3 65400 89800 67000 90000 0 FreeSans 1600 0 0 0 vccd1
port 1 nsew power default
flabel metal3 67400 89800 69000 90000 0 FreeSans 1600 0 0 0 vssd1
port 2 nsew ground default
<< properties >>
string FIXED_BBOX -86 -33820 120052 90020
<< end >>
