magic
tech sky130A
timestamp 1717570567
<< nwell >>
rect -42 133 227 293
rect 427 133 1371 293
<< pwell >>
rect -14 -60 1343 55
<< mvnmos >>
rect 20 0 70 50
rect 99 0 149 50
rect 489 0 539 50
rect 568 0 618 50
rect 706 0 756 50
rect 785 0 835 50
rect 864 0 914 50
rect 943 0 993 50
rect 1022 0 1072 50
rect 1101 0 1151 50
rect 1180 0 1230 50
rect 1259 0 1309 50
<< mvpmos >>
rect 20 166 70 216
rect 99 166 149 216
rect 489 166 539 216
rect 568 166 618 216
rect 706 166 756 216
rect 785 166 835 216
rect 864 166 914 216
rect 943 166 993 216
rect 1022 166 1072 216
rect 1101 166 1151 216
rect 1180 166 1230 216
rect 1259 166 1309 216
<< mvndiff >>
rect -9 46 20 50
rect -9 4 -3 46
rect 14 4 20 46
rect -9 0 20 4
rect 70 46 99 50
rect 70 4 76 46
rect 93 4 99 46
rect 70 0 99 4
rect 149 46 178 50
rect 149 4 155 46
rect 172 4 178 46
rect 149 0 178 4
rect 460 46 489 50
rect 460 4 466 46
rect 483 4 489 46
rect 460 0 489 4
rect 539 46 568 50
rect 539 4 545 46
rect 562 4 568 46
rect 539 0 568 4
rect 618 46 647 50
rect 618 4 624 46
rect 641 4 647 46
rect 618 0 647 4
rect 677 46 706 50
rect 677 4 683 46
rect 700 4 706 46
rect 677 0 706 4
rect 756 46 785 50
rect 756 4 762 46
rect 779 4 785 46
rect 756 0 785 4
rect 835 46 864 50
rect 835 4 841 46
rect 858 4 864 46
rect 835 0 864 4
rect 914 46 943 50
rect 914 4 920 46
rect 937 4 943 46
rect 914 0 943 4
rect 993 46 1022 50
rect 993 4 999 46
rect 1016 4 1022 46
rect 993 0 1022 4
rect 1072 46 1101 50
rect 1072 4 1078 46
rect 1095 4 1101 46
rect 1072 0 1101 4
rect 1151 46 1180 50
rect 1151 4 1157 46
rect 1174 4 1180 46
rect 1151 0 1180 4
rect 1230 46 1259 50
rect 1230 4 1236 46
rect 1253 4 1259 46
rect 1230 0 1259 4
rect 1309 46 1338 50
rect 1309 4 1315 46
rect 1332 4 1338 46
rect 1309 0 1338 4
<< mvpdiff >>
rect -9 212 20 216
rect -9 170 -3 212
rect 14 170 20 212
rect -9 166 20 170
rect 70 212 99 216
rect 70 170 76 212
rect 93 170 99 212
rect 70 166 99 170
rect 149 212 178 216
rect 149 170 155 212
rect 172 170 178 212
rect 149 166 178 170
rect 460 212 489 216
rect 460 170 466 212
rect 483 170 489 212
rect 460 166 489 170
rect 539 212 568 216
rect 539 170 545 212
rect 562 170 568 212
rect 539 166 568 170
rect 618 212 647 216
rect 618 170 624 212
rect 641 170 647 212
rect 618 166 647 170
rect 677 212 706 216
rect 677 170 683 212
rect 700 170 706 212
rect 677 166 706 170
rect 756 212 785 216
rect 756 170 762 212
rect 779 170 785 212
rect 756 166 785 170
rect 835 212 864 216
rect 835 170 841 212
rect 858 170 864 212
rect 835 166 864 170
rect 914 212 943 216
rect 914 170 920 212
rect 937 170 943 212
rect 914 166 943 170
rect 993 212 1022 216
rect 993 170 999 212
rect 1016 170 1022 212
rect 993 166 1022 170
rect 1072 212 1101 216
rect 1072 170 1078 212
rect 1095 170 1101 212
rect 1072 166 1101 170
rect 1151 212 1180 216
rect 1151 170 1157 212
rect 1174 170 1180 212
rect 1151 166 1180 170
rect 1230 212 1259 216
rect 1230 170 1236 212
rect 1253 170 1259 212
rect 1230 166 1259 170
rect 1309 212 1338 216
rect 1309 170 1315 212
rect 1332 170 1338 212
rect 1309 166 1338 170
<< mvndiffc >>
rect -3 4 14 46
rect 76 4 93 46
rect 155 4 172 46
rect 466 4 483 46
rect 545 4 562 46
rect 624 4 641 46
rect 683 4 700 46
rect 762 4 779 46
rect 841 4 858 46
rect 920 4 937 46
rect 999 4 1016 46
rect 1078 4 1095 46
rect 1157 4 1174 46
rect 1236 4 1253 46
rect 1315 4 1332 46
<< mvpdiffc >>
rect -3 170 14 212
rect 76 170 93 212
rect 155 170 172 212
rect 466 170 483 212
rect 545 170 562 212
rect 624 170 641 212
rect 683 170 700 212
rect 762 170 779 212
rect 841 170 858 212
rect 920 170 937 212
rect 999 170 1016 212
rect 1078 170 1095 212
rect 1157 170 1174 212
rect 1236 170 1253 212
rect 1315 170 1332 212
<< mvpsubdiff >>
rect -3 -60 9 -43
rect 1320 -60 1332 -43
<< mvnsubdiff >>
rect -3 243 9 260
rect 182 243 194 260
rect 460 243 472 260
rect 1320 243 1332 260
<< mvpsubdiffcont >>
rect 9 -60 1320 -43
<< mvnsubdiffcont >>
rect 9 243 182 260
rect 472 243 1320 260
<< poly >>
rect 20 216 70 229
rect 99 216 149 229
rect 489 216 539 229
rect 568 216 618 229
rect 706 216 756 229
rect 785 216 835 229
rect 864 216 914 229
rect 943 216 993 229
rect 1022 216 1072 229
rect 1101 216 1151 229
rect 1180 216 1230 229
rect 1259 216 1309 229
rect 20 140 70 166
rect 20 123 31 140
rect 59 123 70 140
rect 20 50 70 123
rect 99 97 149 166
rect 489 142 539 166
rect 489 125 500 142
rect 528 125 539 142
rect 489 120 539 125
rect 568 142 618 166
rect 568 125 579 142
rect 607 125 618 142
rect 568 120 618 125
rect 706 158 756 166
rect 785 158 835 166
rect 864 158 914 166
rect 943 158 993 166
rect 706 131 993 158
rect 99 80 110 97
rect 138 80 149 97
rect 706 114 717 131
rect 745 114 993 131
rect 706 112 993 114
rect 1022 158 1072 166
rect 1101 158 1151 166
rect 1180 158 1230 166
rect 1259 158 1309 166
rect 1022 141 1309 158
rect 99 50 149 80
rect 489 91 539 96
rect 489 74 500 91
rect 528 74 539 91
rect 489 50 539 74
rect 568 91 618 96
rect 568 74 579 91
rect 607 74 618 91
rect 568 50 618 74
rect 706 58 835 112
rect 706 50 756 58
rect 785 50 835 58
rect 864 86 993 91
rect 864 69 880 86
rect 897 69 993 86
rect 864 58 993 69
rect 864 50 914 58
rect 943 50 993 58
rect 1022 75 1027 141
rect 1061 112 1309 141
rect 1061 75 1151 112
rect 1022 58 1151 75
rect 1022 50 1072 58
rect 1101 50 1151 58
rect 1180 86 1309 91
rect 1180 69 1196 86
rect 1213 69 1309 86
rect 1180 58 1309 69
rect 1180 50 1230 58
rect 1259 50 1309 58
rect 20 -13 70 0
rect 99 -13 149 0
rect 489 -13 539 0
rect 568 -13 618 0
rect 706 -13 756 0
rect 785 -13 835 0
rect 864 -13 914 0
rect 943 -13 993 0
rect 1022 -13 1072 0
rect 1101 -13 1151 0
rect 1180 -13 1230 0
rect 1259 -13 1309 0
<< polycont >>
rect 31 123 59 140
rect 500 125 528 142
rect 579 125 607 142
rect 110 80 138 97
rect 717 114 745 131
rect 500 74 528 91
rect 579 74 607 91
rect 880 69 897 86
rect 1027 75 1061 141
rect 1196 69 1213 86
<< locali >>
rect -3 254 9 260
rect 182 254 197 260
rect -3 243 3 254
rect 191 243 197 254
rect 460 254 472 260
rect 1320 254 1332 260
rect 460 243 466 254
rect -3 212 14 220
rect -3 97 14 170
rect 76 212 93 220
rect 76 162 93 170
rect 155 212 172 220
rect 31 140 59 148
rect 31 115 59 123
rect -3 46 14 80
rect 110 97 138 105
rect 110 72 138 80
rect 155 57 172 170
rect -3 -4 14 4
rect 76 46 93 54
rect 76 -21 93 4
rect 155 -4 172 4
rect 466 212 483 220
rect 545 212 562 237
rect 545 162 562 170
rect 624 212 641 220
rect 466 46 483 159
rect 500 142 528 150
rect 500 117 528 125
rect 579 148 584 165
rect 602 148 607 165
rect 579 142 607 148
rect 579 117 607 125
rect 624 139 641 170
rect 683 212 700 237
rect 683 162 700 170
rect 762 212 779 220
rect 762 162 779 170
rect 841 212 858 237
rect 841 162 858 170
rect 920 212 937 220
rect 920 162 937 170
rect 999 212 1016 237
rect 999 162 1016 170
rect 1078 212 1095 220
rect 1027 141 1061 149
rect 624 131 745 139
rect 641 114 717 131
rect 624 106 745 114
rect 500 91 528 99
rect 500 66 528 74
rect 579 91 607 99
rect 579 66 607 74
rect 466 -4 483 4
rect 545 46 562 54
rect 545 -21 562 4
rect 624 46 641 106
rect 841 69 880 86
rect 897 69 937 86
rect 841 54 937 69
rect 1027 67 1061 75
rect 1157 212 1174 237
rect 1157 162 1174 170
rect 1236 212 1253 220
rect 1236 162 1253 170
rect 1315 212 1332 237
rect 1315 162 1332 170
rect 624 -4 641 4
rect 683 46 700 54
rect 683 -21 700 4
rect 762 46 779 54
rect 762 -4 779 4
rect 841 46 858 54
rect 841 -4 858 4
rect 920 46 937 54
rect 920 -4 937 4
rect 999 46 1016 54
rect 999 -4 1016 4
rect 1078 46 1095 132
rect 1078 -4 1095 4
rect 1157 69 1196 86
rect 1213 69 1253 86
rect 1157 54 1253 69
rect 1157 46 1174 54
rect 1157 -4 1174 4
rect 1236 46 1253 54
rect 1236 -4 1253 4
rect 1315 46 1332 54
rect 1315 -4 1332 4
rect 841 -21 1016 -4
rect 1157 -21 1332 -4
rect -3 -43 1332 -38
rect -3 -60 9 -43
rect 1320 -60 1332 -43
<< viali >>
rect 3 243 9 254
rect 9 243 182 254
rect 182 243 191 254
rect 466 243 472 254
rect 472 243 1320 254
rect 1320 243 1332 254
rect 3 237 191 243
rect 466 237 1332 243
rect 76 170 93 212
rect 36 123 54 140
rect -3 80 14 97
rect 115 80 133 97
rect 155 46 172 57
rect 155 40 172 46
rect 466 170 483 176
rect 466 159 483 170
rect 505 125 523 142
rect 584 148 602 165
rect 762 170 779 212
rect 920 170 937 212
rect 1078 170 1095 212
rect 624 114 641 131
rect 722 114 740 131
rect 505 74 523 91
rect 584 74 602 91
rect 1024 75 1027 109
rect 1027 75 1058 109
rect 1078 132 1095 170
rect 1236 170 1253 212
rect 762 4 779 46
rect -3 -38 1332 -21
<< metal1 >>
rect -3 254 197 257
rect -3 237 3 254
rect 191 237 197 254
rect -3 234 197 237
rect 460 254 1338 257
rect 460 237 466 254
rect 1332 237 1338 254
rect 460 234 1338 237
rect 73 212 96 234
rect 762 215 779 218
rect 920 215 937 218
rect 73 170 76 212
rect 93 170 96 212
rect 759 212 782 215
rect 73 164 96 170
rect 463 176 608 182
rect 463 159 466 176
rect 483 165 608 176
rect 759 170 762 212
rect 779 170 782 212
rect 759 167 782 170
rect 917 212 940 215
rect 917 170 920 212
rect 937 170 940 212
rect 917 167 940 170
rect 1075 212 1098 218
rect 1236 215 1253 218
rect 483 159 584 165
rect 463 153 486 159
rect 578 148 584 159
rect 602 148 608 165
rect 30 140 60 148
rect 578 145 608 148
rect 30 123 36 140
rect 54 123 60 140
rect 30 115 60 123
rect 499 142 564 145
rect 499 125 505 142
rect 523 131 564 142
rect 621 134 644 137
rect 621 131 746 134
rect 523 125 624 131
rect 499 122 624 125
rect 543 114 624 122
rect 641 114 722 131
rect 740 114 746 131
rect 621 111 746 114
rect 762 112 779 167
rect 920 112 937 167
rect 1075 132 1078 212
rect 1095 166 1098 212
rect 1233 212 1256 215
rect 1233 170 1236 212
rect 1253 170 1256 212
rect 1233 166 1256 170
rect 1095 132 1371 166
rect 1075 129 1371 132
rect 1078 126 1371 129
rect 621 108 644 111
rect 762 109 1371 112
rect -6 100 17 103
rect -6 97 529 100
rect -6 80 -3 97
rect 14 80 115 97
rect 133 91 529 97
rect 133 80 505 91
rect -6 77 505 80
rect -6 74 17 77
rect 499 74 505 77
rect 523 74 529 91
rect 499 71 529 74
rect 578 91 608 94
rect 578 74 584 91
rect 602 74 608 91
rect 152 57 175 63
rect 578 57 608 74
rect 152 40 155 57
rect 172 40 608 57
rect 762 78 1024 109
rect 762 72 880 78
rect 897 75 1024 78
rect 1058 75 1371 109
rect 897 72 1371 75
rect 762 49 779 72
rect 152 34 608 40
rect 759 46 782 49
rect 759 4 762 46
rect 779 4 782 46
rect 759 1 782 4
rect 762 -2 779 1
rect -9 -21 1338 -18
rect -9 -38 -3 -21
rect 1332 -38 1338 -21
rect -9 -41 1338 -38
<< labels >>
flabel metal1 30 115 60 148 0 FreeSans 160 0 0 0 in
port 1 nsew
flabel locali -3 122 14 139 0 FreeSans 80 90 0 0 in_b
flabel locali 155 116 172 143 0 FreeSans 80 90 0 0 in_bb
flabel metal1 73 234 96 257 0 FreeSans 160 0 0 0 vdd_l
port 4 nsew
flabel metal1 -9 -41 14 -18 0 FreeSans 160 0 0 0 vss
port 6 nsew
flabel metal1 1331 72 1371 112 0 FreeSans 160 0 0 0 out
port 3 nsew
flabel metal1 1331 126 1371 166 0 FreeSans 160 0 0 0 out_b
port 2 nsew
flabel locali 624 80 641 97 0 FreeSans 80 0 0 0 t1
flabel locali 466 116 483 133 0 FreeSans 80 0 0 0 t2
flabel metal1 1315 234 1338 257 0 FreeSans 160 0 0 0 vdd_h
port 5 nsew
<< end >>
