magic
tech sky130A
timestamp 1717520088
<< metal1 >>
rect 3256 44021 3306 44024
rect 3256 43963 3259 44021
rect 3303 43963 3306 44021
rect 3256 41642 3306 43963
rect 16654 44021 16704 44024
rect 16654 43963 16657 44021
rect 16701 43963 16704 44021
rect 3256 41584 3259 41642
rect 3303 41584 3306 41642
rect 3256 41581 3306 41584
rect 3320 43931 3370 43934
rect 3320 43873 3323 43931
rect 3367 43873 3370 43931
rect 3320 41578 3370 43873
rect 16590 43931 16640 43934
rect 16590 43873 16593 43931
rect 16637 43873 16640 43931
rect 3320 41520 3323 41578
rect 3367 41520 3370 41578
rect 3320 41517 3370 41520
rect 3384 42521 3434 42524
rect 3384 42463 3387 42521
rect 3431 42463 3434 42521
rect 3384 41242 3434 42463
rect 16526 42521 16576 42524
rect 16526 42463 16529 42521
rect 16573 42463 16576 42521
rect 3384 41184 3387 41242
rect 3431 41184 3434 41242
rect 3384 41181 3434 41184
rect 3448 42431 3498 42434
rect 3448 42373 3451 42431
rect 3495 42373 3498 42431
rect 3448 41178 3498 42373
rect 16462 42431 16512 42434
rect 16462 42373 16465 42431
rect 16509 42373 16512 42431
rect 3448 41120 3451 41178
rect 3495 41120 3498 41178
rect 3448 41117 3498 41120
rect 3640 41871 5173 41873
rect 3640 41793 5090 41871
rect 5170 41793 5173 41871
rect 14787 41871 16320 41873
rect 14787 41793 14790 41871
rect 14870 41793 16320 41871
rect 3640 41767 3720 41793
rect 5090 41767 5170 41793
rect 3640 41725 5170 41767
rect 3640 41367 3720 41725
rect 3747 41642 3797 41645
rect 3747 41598 3750 41642
rect 3794 41598 3797 41642
rect 3747 41595 3797 41598
rect 4989 41587 5047 41590
rect 3747 41578 3797 41581
rect 3747 41534 3750 41578
rect 3794 41534 3797 41578
rect 3747 41531 3797 41534
rect 4989 41535 4992 41587
rect 5044 41535 5047 41587
rect 4989 41532 5047 41535
rect 5031 41496 5063 41499
rect 5031 41438 5034 41496
rect 5060 41438 5063 41496
rect 5031 41435 5063 41438
rect 5090 41367 5170 41725
rect 14790 41767 14870 41793
rect 16240 41767 16320 41793
rect 14790 41725 16320 41767
rect 3640 41325 5170 41367
rect 3512 41021 3562 41024
rect 3512 40963 3515 41021
rect 3559 40963 3562 41021
rect 3512 40842 3562 40963
rect 3640 40967 3720 41325
rect 3747 41242 3797 41245
rect 3747 41198 3750 41242
rect 3794 41198 3797 41242
rect 3747 41195 3797 41198
rect 4989 41187 5047 41190
rect 3747 41178 3797 41181
rect 3747 41134 3750 41178
rect 3794 41134 3797 41178
rect 3747 41131 3797 41134
rect 4989 41135 4992 41187
rect 5044 41135 5047 41187
rect 4989 41132 5047 41135
rect 5031 41096 5063 41099
rect 5031 41038 5034 41096
rect 5060 41038 5063 41096
rect 5031 41035 5063 41038
rect 5090 41018 5170 41325
rect 14790 41367 14870 41725
rect 16163 41642 16213 41645
rect 16163 41598 16166 41642
rect 16210 41598 16213 41642
rect 16163 41595 16213 41598
rect 14913 41587 14971 41590
rect 14913 41535 14916 41587
rect 14968 41535 14971 41587
rect 14913 41532 14971 41535
rect 16163 41578 16213 41581
rect 16163 41534 16166 41578
rect 16210 41534 16213 41578
rect 16163 41531 16213 41534
rect 14897 41496 14929 41499
rect 14897 41438 14900 41496
rect 14926 41438 14929 41496
rect 14897 41435 14929 41438
rect 16240 41367 16320 41725
rect 14790 41325 16320 41367
rect 14790 41018 14870 41325
rect 16163 41242 16213 41245
rect 16163 41198 16166 41242
rect 16210 41198 16213 41242
rect 16163 41195 16213 41198
rect 14913 41187 14971 41190
rect 14913 41135 14916 41187
rect 14968 41135 14971 41187
rect 14913 41132 14971 41135
rect 16163 41178 16213 41181
rect 16163 41134 16166 41178
rect 16210 41134 16213 41178
rect 16163 41131 16213 41134
rect 14897 41096 14929 41099
rect 14897 41038 14900 41096
rect 14926 41038 14929 41096
rect 14897 41035 14929 41038
rect 5090 40967 5141 41018
rect 3640 40960 5141 40967
rect 5167 40960 5170 41018
rect 14790 40960 14793 41018
rect 14819 40967 14870 41018
rect 16240 40967 16320 41325
rect 16462 41178 16512 42373
rect 16526 41242 16576 42463
rect 16590 41578 16640 43873
rect 16654 41642 16704 43963
rect 16654 41584 16657 41642
rect 16701 41584 16704 41642
rect 16654 41581 16704 41584
rect 16590 41520 16593 41578
rect 16637 41520 16640 41578
rect 16590 41517 16640 41520
rect 16526 41184 16529 41242
rect 16573 41184 16576 41242
rect 16526 41181 16576 41184
rect 16462 41120 16465 41178
rect 16509 41120 16512 41178
rect 16462 41117 16512 41120
rect 14819 40960 16320 40967
rect 3512 40784 3515 40842
rect 3559 40784 3562 40842
rect 3512 40781 3562 40784
rect 3576 40931 3626 40934
rect 3576 40873 3579 40931
rect 3623 40873 3626 40931
rect 3576 40778 3626 40873
rect 3576 40720 3579 40778
rect 3623 40720 3626 40778
rect 3576 40717 3626 40720
rect 3640 40925 5170 40960
rect 3640 40567 3720 40925
rect 3747 40842 3797 40845
rect 3747 40798 3750 40842
rect 3794 40798 3797 40842
rect 3747 40795 3797 40798
rect 4989 40787 5047 40790
rect 3747 40778 3797 40781
rect 3747 40734 3750 40778
rect 3794 40734 3797 40778
rect 3747 40731 3797 40734
rect 4989 40735 4992 40787
rect 5044 40735 5047 40787
rect 4989 40732 5047 40735
rect 5031 40696 5063 40699
rect 5031 40638 5034 40696
rect 5060 40638 5063 40696
rect 5031 40635 5063 40638
rect 5090 40567 5170 40925
rect 14790 40925 16320 40960
rect 16398 41021 16448 41024
rect 16398 40963 16401 41021
rect 16445 40963 16448 41021
rect 3640 40525 5170 40567
rect 3576 40456 3626 40459
rect 3576 40398 3579 40456
rect 3623 40398 3626 40456
rect 3512 40392 3562 40395
rect 3512 40334 3515 40392
rect 3559 40334 3562 40392
rect 3448 40056 3498 40059
rect 3448 39998 3451 40056
rect 3495 39998 3498 40056
rect 3384 39992 3434 39995
rect 3384 39934 3387 39992
rect 3431 39934 3434 39992
rect 3320 39656 3370 39659
rect 3320 39598 3323 39656
rect 3367 39598 3370 39656
rect 3256 39592 3306 39595
rect 3256 39534 3259 39592
rect 3303 39534 3306 39592
rect 3192 39256 3242 39259
rect 3192 39198 3195 39256
rect 3239 39198 3242 39256
rect 3128 39192 3178 39195
rect 3128 39134 3131 39192
rect 3175 39134 3178 39192
rect 3064 38856 3114 38859
rect 3064 38798 3067 38856
rect 3111 38798 3114 38856
rect 3000 38792 3050 38795
rect 3000 38734 3003 38792
rect 3047 38734 3050 38792
rect 2936 38456 2986 38459
rect 2936 38398 2939 38456
rect 2983 38398 2986 38456
rect 2872 38392 2922 38395
rect 2872 38334 2875 38392
rect 2919 38334 2922 38392
rect 2808 38155 2858 38158
rect 2808 38097 2811 38155
rect 2855 38097 2858 38155
rect 2744 38091 2794 38094
rect 2744 38033 2747 38091
rect 2791 38033 2794 38091
rect 2680 37656 2730 37659
rect 2680 37598 2683 37656
rect 2727 37598 2730 37656
rect 2616 37592 2666 37595
rect 2616 37534 2619 37592
rect 2663 37534 2666 37592
rect 2552 37256 2602 37259
rect 2552 37198 2555 37256
rect 2599 37198 2602 37256
rect 2488 37192 2538 37195
rect 2488 37134 2491 37192
rect 2535 37134 2538 37192
rect 2424 36856 2474 36859
rect 2424 36798 2427 36856
rect 2471 36798 2474 36856
rect 2360 36792 2410 36795
rect 2360 36734 2363 36792
rect 2407 36734 2410 36792
rect 2296 36655 2346 36658
rect 2296 36597 2299 36655
rect 2343 36597 2346 36655
rect 2232 36591 2282 36594
rect 2232 36533 2235 36591
rect 2279 36533 2282 36591
rect 2168 36056 2218 36059
rect 2168 35998 2171 36056
rect 2215 35998 2218 36056
rect 2104 35992 2154 35995
rect 2104 35934 2107 35992
rect 2151 35934 2154 35992
rect 2040 35656 2090 35659
rect 2040 35598 2043 35656
rect 2087 35598 2090 35656
rect 1976 35592 2026 35595
rect 1976 35534 1979 35592
rect 2023 35534 2026 35592
rect 1912 35256 1962 35259
rect 1912 35198 1915 35256
rect 1959 35198 1962 35256
rect 1848 35192 1898 35195
rect 1848 35134 1851 35192
rect 1895 35134 1898 35192
rect 1784 34853 1834 34856
rect 1784 34795 1787 34853
rect 1831 34795 1834 34853
rect 1720 34789 1770 34792
rect 1720 34731 1723 34789
rect 1767 34731 1770 34789
rect 1656 34456 1706 34459
rect 1656 34398 1659 34456
rect 1703 34398 1706 34456
rect 1592 34392 1642 34395
rect 1592 34334 1595 34392
rect 1639 34334 1642 34392
rect 1528 34056 1578 34059
rect 1528 33998 1531 34056
rect 1575 33998 1578 34056
rect 1464 33992 1514 33995
rect 1464 33934 1467 33992
rect 1511 33934 1514 33992
rect 1400 33656 1450 33659
rect 1400 33598 1403 33656
rect 1447 33598 1450 33656
rect 1336 33592 1386 33595
rect 1336 33534 1339 33592
rect 1383 33534 1386 33592
rect 1272 33256 1322 33259
rect 1272 33198 1275 33256
rect 1319 33198 1322 33256
rect 1208 33192 1258 33195
rect 1208 33134 1211 33192
rect 1255 33134 1258 33192
rect 1144 32856 1194 32859
rect 1144 32798 1147 32856
rect 1191 32798 1194 32856
rect 1080 32792 1130 32795
rect 1080 32734 1083 32792
rect 1127 32734 1130 32792
rect 1016 32456 1066 32459
rect 1016 32398 1019 32456
rect 1063 32398 1066 32456
rect 952 32392 1002 32395
rect 952 32334 955 32392
rect 999 32334 1002 32392
rect 888 32149 938 32152
rect 888 32091 891 32149
rect 935 32091 938 32149
rect 824 32085 874 32088
rect 824 32027 827 32085
rect 871 32027 874 32085
rect 760 31656 810 31659
rect 760 31598 763 31656
rect 807 31598 810 31656
rect 696 31592 746 31595
rect 696 31534 699 31592
rect 743 31534 746 31592
rect 632 31256 682 31259
rect 632 31198 635 31256
rect 679 31198 682 31256
rect 568 31192 618 31195
rect 568 31134 571 31192
rect 615 31134 618 31192
rect 504 30856 554 30859
rect 504 30798 507 30856
rect 551 30798 554 30856
rect 440 30792 490 30795
rect 440 30734 443 30792
rect 487 30734 490 30792
rect 376 30655 426 30658
rect 376 30597 379 30655
rect 423 30597 426 30655
rect 312 30591 362 30594
rect 312 30533 315 30591
rect 359 30533 362 30591
rect 248 30056 298 30059
rect 248 29998 251 30056
rect 295 29998 298 30056
rect 184 29992 234 29995
rect 184 29934 187 29992
rect 231 29934 234 29992
rect 184 417 234 29934
rect 248 507 298 29998
rect 312 1917 362 30533
rect 376 2007 426 30597
rect 440 3417 490 30734
rect 504 3507 554 30798
rect 568 4917 618 31134
rect 632 5007 682 31198
rect 696 6417 746 31534
rect 760 6507 810 31598
rect 824 7917 874 32027
rect 888 8007 938 32091
rect 952 9417 1002 32334
rect 1016 9507 1066 32398
rect 1080 10917 1130 32734
rect 1144 11007 1194 32798
rect 1208 12417 1258 33134
rect 1272 12507 1322 33198
rect 1336 13917 1386 33534
rect 1400 14007 1450 33598
rect 1464 15417 1514 33934
rect 1528 15507 1578 33998
rect 1592 16917 1642 34334
rect 1656 17007 1706 34398
rect 1720 18417 1770 34731
rect 1784 18507 1834 34795
rect 1848 19917 1898 35134
rect 1912 20007 1962 35198
rect 1976 21417 2026 35534
rect 2040 21507 2090 35598
rect 2104 22917 2154 35934
rect 2168 23007 2218 35998
rect 2232 24417 2282 36533
rect 2296 24507 2346 36597
rect 2360 25917 2410 36734
rect 2424 26007 2474 36798
rect 2488 27417 2538 37134
rect 2552 27507 2602 37198
rect 2616 28917 2666 37534
rect 2680 29007 2730 37598
rect 2744 30417 2794 38033
rect 2808 30507 2858 38097
rect 2872 31917 2922 38334
rect 2936 32007 2986 38398
rect 3000 33417 3050 38734
rect 3064 33507 3114 38798
rect 3128 34917 3178 39134
rect 3192 35007 3242 39198
rect 3256 36417 3306 39534
rect 3320 36507 3370 39598
rect 3384 37917 3434 39934
rect 3448 38007 3498 39998
rect 3512 39417 3562 40334
rect 3576 39507 3626 40398
rect 3576 39449 3579 39507
rect 3623 39449 3626 39507
rect 3576 39446 3626 39449
rect 3640 40167 3720 40525
rect 3747 40442 3797 40445
rect 3747 40398 3750 40442
rect 3794 40398 3797 40442
rect 3747 40395 3797 40398
rect 4989 40387 5047 40390
rect 3747 40378 3797 40381
rect 3747 40334 3750 40378
rect 3794 40334 3797 40378
rect 3747 40331 3797 40334
rect 4989 40335 4992 40387
rect 5044 40335 5047 40387
rect 4989 40332 5047 40335
rect 5031 40296 5063 40299
rect 5031 40238 5034 40296
rect 5060 40238 5063 40296
rect 5031 40235 5063 40238
rect 5090 40218 5170 40525
rect 14790 40567 14870 40925
rect 16163 40842 16213 40845
rect 16163 40798 16166 40842
rect 16210 40798 16213 40842
rect 16163 40795 16213 40798
rect 14913 40787 14971 40790
rect 14913 40735 14916 40787
rect 14968 40735 14971 40787
rect 14913 40732 14971 40735
rect 16163 40778 16213 40781
rect 16163 40734 16166 40778
rect 16210 40734 16213 40778
rect 16163 40731 16213 40734
rect 14897 40696 14929 40699
rect 14897 40638 14900 40696
rect 14926 40638 14929 40696
rect 14897 40635 14929 40638
rect 16240 40567 16320 40925
rect 16334 40931 16384 40934
rect 16334 40873 16337 40931
rect 16381 40873 16384 40931
rect 16334 40778 16384 40873
rect 16398 40842 16448 40963
rect 16398 40784 16401 40842
rect 16445 40784 16448 40842
rect 16398 40781 16448 40784
rect 16334 40720 16337 40778
rect 16381 40720 16384 40778
rect 16334 40717 16384 40720
rect 14790 40525 16320 40567
rect 14790 40218 14870 40525
rect 16163 40442 16213 40445
rect 16163 40398 16166 40442
rect 16210 40398 16213 40442
rect 16163 40395 16213 40398
rect 14913 40387 14971 40390
rect 14913 40335 14916 40387
rect 14968 40335 14971 40387
rect 14913 40332 14971 40335
rect 16163 40378 16213 40381
rect 16163 40334 16166 40378
rect 16210 40334 16213 40378
rect 16163 40331 16213 40334
rect 14897 40296 14929 40299
rect 14897 40238 14900 40296
rect 14926 40238 14929 40296
rect 14897 40235 14929 40238
rect 5090 40167 5141 40218
rect 3640 40160 5141 40167
rect 5167 40160 5170 40218
rect 14790 40160 14793 40218
rect 14819 40167 14870 40218
rect 16240 40167 16320 40525
rect 14819 40160 16320 40167
rect 3640 40125 5170 40160
rect 3640 39767 3720 40125
rect 3747 40042 3797 40045
rect 3747 39998 3750 40042
rect 3794 39998 3797 40042
rect 3747 39995 3797 39998
rect 4989 39987 5047 39990
rect 3747 39978 3797 39981
rect 3747 39934 3750 39978
rect 3794 39934 3797 39978
rect 3747 39931 3797 39934
rect 4989 39935 4992 39987
rect 5044 39935 5047 39987
rect 4989 39932 5047 39935
rect 5031 39896 5063 39899
rect 5031 39838 5034 39896
rect 5060 39838 5063 39896
rect 5031 39835 5063 39838
rect 5090 39767 5170 40125
rect 14790 40125 16320 40160
rect 3640 39725 5170 39767
rect 3512 39359 3515 39417
rect 3559 39359 3562 39417
rect 3512 39356 3562 39359
rect 3640 39367 3720 39725
rect 3747 39642 3797 39645
rect 3747 39598 3750 39642
rect 3794 39598 3797 39642
rect 3747 39595 3797 39598
rect 4989 39587 5047 39590
rect 3747 39578 3797 39581
rect 3747 39534 3750 39578
rect 3794 39534 3797 39578
rect 3747 39531 3797 39534
rect 4989 39535 4992 39587
rect 5044 39535 5047 39587
rect 4989 39532 5047 39535
rect 5031 39496 5063 39499
rect 5031 39438 5034 39496
rect 5060 39438 5063 39496
rect 5031 39435 5063 39438
rect 5090 39418 5170 39725
rect 14790 39767 14870 40125
rect 16163 40042 16213 40045
rect 16163 39998 16166 40042
rect 16210 39998 16213 40042
rect 16163 39995 16213 39998
rect 14913 39987 14971 39990
rect 14913 39935 14916 39987
rect 14968 39935 14971 39987
rect 14913 39932 14971 39935
rect 16163 39978 16213 39981
rect 16163 39934 16166 39978
rect 16210 39934 16213 39978
rect 16163 39931 16213 39934
rect 14897 39896 14929 39899
rect 14897 39838 14900 39896
rect 14926 39838 14929 39896
rect 14897 39835 14929 39838
rect 16240 39767 16320 40125
rect 14790 39725 16320 39767
rect 14790 39418 14870 39725
rect 16163 39642 16213 39645
rect 16163 39598 16166 39642
rect 16210 39598 16213 39642
rect 16163 39595 16213 39598
rect 14913 39587 14971 39590
rect 14913 39535 14916 39587
rect 14968 39535 14971 39587
rect 14913 39532 14971 39535
rect 16163 39578 16213 39581
rect 16163 39534 16166 39578
rect 16210 39534 16213 39578
rect 16163 39531 16213 39534
rect 14897 39496 14929 39499
rect 14897 39438 14900 39496
rect 14926 39438 14929 39496
rect 14897 39435 14929 39438
rect 5090 39367 5141 39418
rect 3640 39360 5141 39367
rect 5167 39360 5170 39418
rect 14790 39360 14793 39418
rect 14819 39367 14870 39418
rect 16240 39367 16320 39725
rect 16334 40456 16384 40459
rect 16334 40398 16337 40456
rect 16381 40398 16384 40456
rect 16334 39507 16384 40398
rect 16334 39449 16337 39507
rect 16381 39449 16384 39507
rect 16334 39446 16384 39449
rect 16398 40392 16448 40395
rect 16398 40334 16401 40392
rect 16445 40334 16448 40392
rect 14819 39360 16320 39367
rect 3448 37949 3451 38007
rect 3495 37949 3498 38007
rect 3448 37946 3498 37949
rect 3640 39325 5170 39360
rect 3640 38967 3720 39325
rect 3747 39242 3797 39245
rect 3747 39198 3750 39242
rect 3794 39198 3797 39242
rect 3747 39195 3797 39198
rect 4989 39187 5047 39190
rect 3747 39178 3797 39181
rect 3747 39134 3750 39178
rect 3794 39134 3797 39178
rect 3747 39131 3797 39134
rect 4989 39135 4992 39187
rect 5044 39135 5047 39187
rect 4989 39132 5047 39135
rect 5031 39096 5063 39099
rect 5031 39038 5034 39096
rect 5060 39038 5063 39096
rect 5031 39035 5063 39038
rect 5090 38967 5170 39325
rect 14790 39325 16320 39360
rect 16398 39417 16448 40334
rect 16398 39359 16401 39417
rect 16445 39359 16448 39417
rect 16398 39356 16448 39359
rect 16462 40056 16512 40059
rect 16462 39998 16465 40056
rect 16509 39998 16512 40056
rect 3640 38925 5170 38967
rect 3640 38567 3720 38925
rect 3747 38842 3797 38845
rect 3747 38798 3750 38842
rect 3794 38798 3797 38842
rect 3747 38795 3797 38798
rect 4989 38787 5047 38790
rect 3747 38778 3797 38781
rect 3747 38734 3750 38778
rect 3794 38734 3797 38778
rect 3747 38731 3797 38734
rect 4989 38735 4992 38787
rect 5044 38735 5047 38787
rect 4989 38732 5047 38735
rect 5031 38696 5063 38699
rect 5031 38638 5034 38696
rect 5060 38638 5063 38696
rect 5031 38635 5063 38638
rect 5090 38618 5170 38925
rect 14790 38967 14870 39325
rect 16163 39242 16213 39245
rect 16163 39198 16166 39242
rect 16210 39198 16213 39242
rect 16163 39195 16213 39198
rect 14913 39187 14971 39190
rect 14913 39135 14916 39187
rect 14968 39135 14971 39187
rect 14913 39132 14971 39135
rect 16163 39178 16213 39181
rect 16163 39134 16166 39178
rect 16210 39134 16213 39178
rect 16163 39131 16213 39134
rect 14897 39096 14929 39099
rect 14897 39038 14900 39096
rect 14926 39038 14929 39096
rect 14897 39035 14929 39038
rect 16240 38967 16320 39325
rect 14790 38925 16320 38967
rect 14790 38618 14870 38925
rect 16163 38842 16213 38845
rect 16163 38798 16166 38842
rect 16210 38798 16213 38842
rect 16163 38795 16213 38798
rect 14913 38787 14971 38790
rect 14913 38735 14916 38787
rect 14968 38735 14971 38787
rect 14913 38732 14971 38735
rect 16163 38778 16213 38781
rect 16163 38734 16166 38778
rect 16210 38734 16213 38778
rect 16163 38731 16213 38734
rect 14897 38696 14929 38699
rect 14897 38638 14900 38696
rect 14926 38638 14929 38696
rect 14897 38635 14929 38638
rect 5090 38567 5141 38618
rect 3640 38560 5141 38567
rect 5167 38560 5170 38618
rect 14790 38560 14793 38618
rect 14819 38567 14870 38618
rect 16240 38567 16320 38925
rect 14819 38560 16320 38567
rect 3640 38525 5170 38560
rect 3640 38167 3720 38525
rect 3747 38442 3797 38445
rect 3747 38398 3750 38442
rect 3794 38398 3797 38442
rect 3747 38395 3797 38398
rect 4989 38387 5047 38390
rect 3747 38378 3797 38381
rect 3747 38334 3750 38378
rect 3794 38334 3797 38378
rect 3747 38331 3797 38334
rect 4989 38335 4992 38387
rect 5044 38335 5047 38387
rect 4989 38332 5047 38335
rect 5031 38296 5063 38299
rect 5031 38238 5034 38296
rect 5060 38238 5063 38296
rect 5031 38235 5063 38238
rect 5090 38167 5170 38525
rect 14790 38525 16320 38560
rect 3640 38125 5170 38167
rect 3384 37859 3387 37917
rect 3431 37859 3434 37917
rect 3384 37856 3434 37859
rect 3320 36449 3323 36507
rect 3367 36449 3370 36507
rect 3320 36446 3370 36449
rect 3640 37767 3720 38125
rect 3747 38042 3797 38045
rect 3747 37998 3750 38042
rect 3794 37998 3797 38042
rect 3747 37995 3797 37998
rect 4989 37987 5047 37990
rect 3747 37978 3797 37981
rect 3747 37934 3750 37978
rect 3794 37934 3797 37978
rect 3747 37931 3797 37934
rect 4989 37935 4992 37987
rect 5044 37935 5047 37987
rect 4989 37932 5047 37935
rect 5031 37896 5063 37899
rect 5031 37838 5034 37896
rect 5060 37838 5063 37896
rect 5031 37835 5063 37838
rect 5090 37818 5170 38125
rect 14790 38167 14870 38525
rect 16163 38442 16213 38445
rect 16163 38398 16166 38442
rect 16210 38398 16213 38442
rect 16163 38395 16213 38398
rect 14913 38387 14971 38390
rect 14913 38335 14916 38387
rect 14968 38335 14971 38387
rect 14913 38332 14971 38335
rect 16163 38378 16213 38381
rect 16163 38334 16166 38378
rect 16210 38334 16213 38378
rect 16163 38331 16213 38334
rect 14897 38296 14929 38299
rect 14897 38238 14900 38296
rect 14926 38238 14929 38296
rect 14897 38235 14929 38238
rect 16240 38167 16320 38525
rect 14790 38125 16320 38167
rect 14790 37818 14870 38125
rect 16163 38042 16213 38045
rect 16163 37998 16166 38042
rect 16210 37998 16213 38042
rect 16163 37995 16213 37998
rect 14913 37987 14971 37990
rect 14913 37935 14916 37987
rect 14968 37935 14971 37987
rect 14913 37932 14971 37935
rect 16163 37978 16213 37981
rect 16163 37934 16166 37978
rect 16210 37934 16213 37978
rect 16163 37931 16213 37934
rect 14897 37896 14929 37899
rect 14897 37838 14900 37896
rect 14926 37838 14929 37896
rect 14897 37835 14929 37838
rect 5090 37767 5141 37818
rect 3640 37760 5141 37767
rect 5167 37760 5170 37818
rect 14790 37760 14793 37818
rect 14819 37767 14870 37818
rect 16240 37767 16320 38125
rect 16462 38007 16512 39998
rect 16462 37949 16465 38007
rect 16509 37949 16512 38007
rect 16462 37946 16512 37949
rect 16526 39992 16576 39995
rect 16526 39934 16529 39992
rect 16573 39934 16576 39992
rect 16526 37917 16576 39934
rect 16526 37859 16529 37917
rect 16573 37859 16576 37917
rect 16526 37856 16576 37859
rect 16590 39656 16640 39659
rect 16590 39598 16593 39656
rect 16637 39598 16640 39656
rect 14819 37760 16320 37767
rect 3640 37725 5170 37760
rect 3640 37367 3720 37725
rect 3747 37642 3797 37645
rect 3747 37598 3750 37642
rect 3794 37598 3797 37642
rect 3747 37595 3797 37598
rect 4989 37587 5047 37590
rect 3747 37578 3797 37581
rect 3747 37534 3750 37578
rect 3794 37534 3797 37578
rect 3747 37531 3797 37534
rect 4989 37535 4992 37587
rect 5044 37535 5047 37587
rect 4989 37532 5047 37535
rect 5031 37496 5063 37499
rect 5031 37438 5034 37496
rect 5060 37438 5063 37496
rect 5031 37435 5063 37438
rect 5090 37367 5170 37725
rect 14790 37725 16320 37760
rect 3640 37325 5170 37367
rect 3640 36967 3720 37325
rect 3747 37242 3797 37245
rect 3747 37198 3750 37242
rect 3794 37198 3797 37242
rect 3747 37195 3797 37198
rect 4989 37187 5047 37190
rect 3747 37178 3797 37181
rect 3747 37134 3750 37178
rect 3794 37134 3797 37178
rect 3747 37131 3797 37134
rect 4989 37135 4992 37187
rect 5044 37135 5047 37187
rect 4989 37132 5047 37135
rect 5031 37096 5063 37099
rect 5031 37038 5034 37096
rect 5060 37038 5063 37096
rect 5031 37035 5063 37038
rect 5090 37018 5170 37325
rect 14790 37367 14870 37725
rect 16163 37642 16213 37645
rect 16163 37598 16166 37642
rect 16210 37598 16213 37642
rect 16163 37595 16213 37598
rect 14913 37587 14971 37590
rect 14913 37535 14916 37587
rect 14968 37535 14971 37587
rect 14913 37532 14971 37535
rect 16163 37578 16213 37581
rect 16163 37534 16166 37578
rect 16210 37534 16213 37578
rect 16163 37531 16213 37534
rect 14897 37496 14929 37499
rect 14897 37438 14900 37496
rect 14926 37438 14929 37496
rect 14897 37435 14929 37438
rect 16240 37367 16320 37725
rect 14790 37325 16320 37367
rect 14790 37018 14870 37325
rect 16163 37242 16213 37245
rect 16163 37198 16166 37242
rect 16210 37198 16213 37242
rect 16163 37195 16213 37198
rect 14913 37187 14971 37190
rect 14913 37135 14916 37187
rect 14968 37135 14971 37187
rect 14913 37132 14971 37135
rect 16163 37178 16213 37181
rect 16163 37134 16166 37178
rect 16210 37134 16213 37178
rect 16163 37131 16213 37134
rect 14897 37096 14929 37099
rect 14897 37038 14900 37096
rect 14926 37038 14929 37096
rect 14897 37035 14929 37038
rect 5090 36967 5141 37018
rect 3640 36960 5141 36967
rect 5167 36960 5170 37018
rect 14790 36960 14793 37018
rect 14819 36967 14870 37018
rect 16240 36967 16320 37325
rect 14819 36960 16320 36967
rect 3640 36925 5170 36960
rect 3640 36567 3720 36925
rect 3747 36842 3797 36845
rect 3747 36798 3750 36842
rect 3794 36798 3797 36842
rect 3747 36795 3797 36798
rect 4989 36787 5047 36790
rect 3747 36778 3797 36781
rect 3747 36734 3750 36778
rect 3794 36734 3797 36778
rect 3747 36731 3797 36734
rect 4989 36735 4992 36787
rect 5044 36735 5047 36787
rect 4989 36732 5047 36735
rect 5031 36696 5063 36699
rect 5031 36638 5034 36696
rect 5060 36638 5063 36696
rect 5031 36635 5063 36638
rect 5090 36567 5170 36925
rect 14790 36925 16320 36960
rect 3640 36525 5170 36567
rect 3256 36359 3259 36417
rect 3303 36359 3306 36417
rect 3256 36356 3306 36359
rect 3192 34949 3195 35007
rect 3239 34949 3242 35007
rect 3192 34946 3242 34949
rect 3640 36167 3720 36525
rect 3747 36442 3797 36445
rect 3747 36398 3750 36442
rect 3794 36398 3797 36442
rect 3747 36395 3797 36398
rect 4989 36387 5047 36390
rect 3747 36378 3797 36381
rect 3747 36334 3750 36378
rect 3794 36334 3797 36378
rect 3747 36331 3797 36334
rect 4989 36335 4992 36387
rect 5044 36335 5047 36387
rect 4989 36332 5047 36335
rect 5031 36296 5063 36299
rect 5031 36238 5034 36296
rect 5060 36238 5063 36296
rect 5031 36235 5063 36238
rect 5090 36218 5170 36525
rect 14790 36567 14870 36925
rect 16163 36842 16213 36845
rect 16163 36798 16166 36842
rect 16210 36798 16213 36842
rect 16163 36795 16213 36798
rect 14913 36787 14971 36790
rect 14913 36735 14916 36787
rect 14968 36735 14971 36787
rect 14913 36732 14971 36735
rect 16163 36778 16213 36781
rect 16163 36734 16166 36778
rect 16210 36734 16213 36778
rect 16163 36731 16213 36734
rect 14897 36696 14929 36699
rect 14897 36638 14900 36696
rect 14926 36638 14929 36696
rect 14897 36635 14929 36638
rect 16240 36567 16320 36925
rect 14790 36525 16320 36567
rect 14790 36218 14870 36525
rect 16163 36442 16213 36445
rect 16163 36398 16166 36442
rect 16210 36398 16213 36442
rect 16163 36395 16213 36398
rect 14913 36387 14971 36390
rect 14913 36335 14916 36387
rect 14968 36335 14971 36387
rect 14913 36332 14971 36335
rect 16163 36378 16213 36381
rect 16163 36334 16166 36378
rect 16210 36334 16213 36378
rect 16163 36331 16213 36334
rect 14897 36296 14929 36299
rect 14897 36238 14900 36296
rect 14926 36238 14929 36296
rect 14897 36235 14929 36238
rect 5090 36167 5141 36218
rect 3640 36160 5141 36167
rect 5167 36160 5170 36218
rect 14790 36160 14793 36218
rect 14819 36167 14870 36218
rect 16240 36167 16320 36525
rect 16590 36507 16640 39598
rect 16590 36449 16593 36507
rect 16637 36449 16640 36507
rect 16590 36446 16640 36449
rect 16654 39592 16704 39595
rect 16654 39534 16657 39592
rect 16701 39534 16704 39592
rect 16654 36417 16704 39534
rect 16654 36359 16657 36417
rect 16701 36359 16704 36417
rect 16654 36356 16704 36359
rect 16718 39256 16768 39259
rect 16718 39198 16721 39256
rect 16765 39198 16768 39256
rect 14819 36160 16320 36167
rect 3640 36125 5170 36160
rect 3640 35767 3720 36125
rect 3747 36042 3797 36045
rect 3747 35998 3750 36042
rect 3794 35998 3797 36042
rect 3747 35995 3797 35998
rect 4989 35987 5047 35990
rect 3747 35978 3797 35981
rect 3747 35934 3750 35978
rect 3794 35934 3797 35978
rect 3747 35931 3797 35934
rect 4989 35935 4992 35987
rect 5044 35935 5047 35987
rect 4989 35932 5047 35935
rect 5031 35896 5063 35899
rect 5031 35838 5034 35896
rect 5060 35838 5063 35896
rect 5031 35835 5063 35838
rect 5090 35767 5170 36125
rect 14790 36125 16320 36160
rect 3640 35725 5170 35767
rect 3640 35367 3720 35725
rect 3747 35642 3797 35645
rect 3747 35598 3750 35642
rect 3794 35598 3797 35642
rect 3747 35595 3797 35598
rect 4989 35587 5047 35590
rect 3747 35578 3797 35581
rect 3747 35534 3750 35578
rect 3794 35534 3797 35578
rect 3747 35531 3797 35534
rect 4989 35535 4992 35587
rect 5044 35535 5047 35587
rect 4989 35532 5047 35535
rect 5031 35496 5063 35499
rect 5031 35438 5034 35496
rect 5060 35438 5063 35496
rect 5031 35435 5063 35438
rect 5090 35418 5170 35725
rect 14790 35767 14870 36125
rect 16163 36042 16213 36045
rect 16163 35998 16166 36042
rect 16210 35998 16213 36042
rect 16163 35995 16213 35998
rect 14913 35987 14971 35990
rect 14913 35935 14916 35987
rect 14968 35935 14971 35987
rect 14913 35932 14971 35935
rect 16163 35978 16213 35981
rect 16163 35934 16166 35978
rect 16210 35934 16213 35978
rect 16163 35931 16213 35934
rect 14897 35896 14929 35899
rect 14897 35838 14900 35896
rect 14926 35838 14929 35896
rect 14897 35835 14929 35838
rect 16240 35767 16320 36125
rect 14790 35725 16320 35767
rect 14790 35418 14870 35725
rect 16163 35642 16213 35645
rect 16163 35598 16166 35642
rect 16210 35598 16213 35642
rect 16163 35595 16213 35598
rect 14913 35587 14971 35590
rect 14913 35535 14916 35587
rect 14968 35535 14971 35587
rect 14913 35532 14971 35535
rect 16163 35578 16213 35581
rect 16163 35534 16166 35578
rect 16210 35534 16213 35578
rect 16163 35531 16213 35534
rect 14897 35496 14929 35499
rect 14897 35438 14900 35496
rect 14926 35438 14929 35496
rect 14897 35435 14929 35438
rect 5090 35367 5141 35418
rect 3640 35360 5141 35367
rect 5167 35360 5170 35418
rect 14790 35360 14793 35418
rect 14819 35367 14870 35418
rect 16240 35367 16320 35725
rect 14819 35360 16320 35367
rect 3640 35325 5170 35360
rect 3640 34967 3720 35325
rect 3747 35242 3797 35245
rect 3747 35198 3750 35242
rect 3794 35198 3797 35242
rect 3747 35195 3797 35198
rect 4989 35187 5047 35190
rect 3747 35178 3797 35181
rect 3747 35134 3750 35178
rect 3794 35134 3797 35178
rect 3747 35131 3797 35134
rect 4989 35135 4992 35187
rect 5044 35135 5047 35187
rect 4989 35132 5047 35135
rect 5031 35096 5063 35099
rect 5031 35038 5034 35096
rect 5060 35038 5063 35096
rect 5031 35035 5063 35038
rect 5090 34967 5170 35325
rect 14790 35325 16320 35360
rect 3128 34859 3131 34917
rect 3175 34859 3178 34917
rect 3128 34856 3178 34859
rect 3640 34925 5170 34967
rect 3064 33449 3067 33507
rect 3111 33449 3114 33507
rect 3064 33446 3114 33449
rect 3640 34567 3720 34925
rect 3747 34842 3797 34845
rect 3747 34798 3750 34842
rect 3794 34798 3797 34842
rect 3747 34795 3797 34798
rect 4989 34787 5047 34790
rect 3747 34778 3797 34781
rect 3747 34734 3750 34778
rect 3794 34734 3797 34778
rect 3747 34731 3797 34734
rect 4989 34735 4992 34787
rect 5044 34735 5047 34787
rect 4989 34732 5047 34735
rect 5031 34696 5063 34699
rect 5031 34638 5034 34696
rect 5060 34638 5063 34696
rect 5031 34635 5063 34638
rect 5090 34618 5170 34925
rect 14790 34967 14870 35325
rect 16163 35242 16213 35245
rect 16163 35198 16166 35242
rect 16210 35198 16213 35242
rect 16163 35195 16213 35198
rect 14913 35187 14971 35190
rect 14913 35135 14916 35187
rect 14968 35135 14971 35187
rect 14913 35132 14971 35135
rect 16163 35178 16213 35181
rect 16163 35134 16166 35178
rect 16210 35134 16213 35178
rect 16163 35131 16213 35134
rect 14897 35096 14929 35099
rect 14897 35038 14900 35096
rect 14926 35038 14929 35096
rect 14897 35035 14929 35038
rect 16240 34967 16320 35325
rect 14790 34925 16320 34967
rect 16718 35007 16768 39198
rect 16718 34949 16721 35007
rect 16765 34949 16768 35007
rect 16718 34946 16768 34949
rect 16782 39192 16832 39195
rect 16782 39134 16785 39192
rect 16829 39134 16832 39192
rect 14790 34618 14870 34925
rect 16163 34842 16213 34845
rect 16163 34798 16166 34842
rect 16210 34798 16213 34842
rect 16163 34795 16213 34798
rect 14913 34787 14971 34790
rect 14913 34735 14916 34787
rect 14968 34735 14971 34787
rect 14913 34732 14971 34735
rect 16163 34778 16213 34781
rect 16163 34734 16166 34778
rect 16210 34734 16213 34778
rect 16163 34731 16213 34734
rect 14897 34696 14929 34699
rect 14897 34638 14900 34696
rect 14926 34638 14929 34696
rect 14897 34635 14929 34638
rect 5090 34567 5141 34618
rect 3640 34560 5141 34567
rect 5167 34560 5170 34618
rect 14790 34560 14793 34618
rect 14819 34567 14870 34618
rect 16240 34567 16320 34925
rect 16782 34917 16832 39134
rect 16782 34859 16785 34917
rect 16829 34859 16832 34917
rect 16782 34856 16832 34859
rect 16846 38856 16896 38859
rect 16846 38798 16849 38856
rect 16893 38798 16896 38856
rect 14819 34560 16320 34567
rect 3640 34525 5170 34560
rect 3640 34167 3720 34525
rect 3747 34442 3797 34445
rect 3747 34398 3750 34442
rect 3794 34398 3797 34442
rect 3747 34395 3797 34398
rect 4989 34387 5047 34390
rect 3747 34378 3797 34381
rect 3747 34334 3750 34378
rect 3794 34334 3797 34378
rect 3747 34331 3797 34334
rect 4989 34335 4992 34387
rect 5044 34335 5047 34387
rect 4989 34332 5047 34335
rect 5031 34296 5063 34299
rect 5031 34238 5034 34296
rect 5060 34238 5063 34296
rect 5031 34235 5063 34238
rect 5090 34167 5170 34525
rect 14790 34525 16320 34560
rect 3640 34125 5170 34167
rect 3640 33767 3720 34125
rect 3747 34042 3797 34045
rect 3747 33998 3750 34042
rect 3794 33998 3797 34042
rect 3747 33995 3797 33998
rect 4989 33987 5047 33990
rect 3747 33978 3797 33981
rect 3747 33934 3750 33978
rect 3794 33934 3797 33978
rect 3747 33931 3797 33934
rect 4989 33935 4992 33987
rect 5044 33935 5047 33987
rect 4989 33932 5047 33935
rect 5031 33896 5063 33899
rect 5031 33838 5034 33896
rect 5060 33838 5063 33896
rect 5031 33835 5063 33838
rect 5090 33818 5170 34125
rect 14790 34167 14870 34525
rect 16163 34442 16213 34445
rect 16163 34398 16166 34442
rect 16210 34398 16213 34442
rect 16163 34395 16213 34398
rect 14913 34387 14971 34390
rect 14913 34335 14916 34387
rect 14968 34335 14971 34387
rect 14913 34332 14971 34335
rect 16163 34378 16213 34381
rect 16163 34334 16166 34378
rect 16210 34334 16213 34378
rect 16163 34331 16213 34334
rect 14897 34296 14929 34299
rect 14897 34238 14900 34296
rect 14926 34238 14929 34296
rect 14897 34235 14929 34238
rect 16240 34167 16320 34525
rect 14790 34125 16320 34167
rect 14790 33818 14870 34125
rect 16163 34042 16213 34045
rect 16163 33998 16166 34042
rect 16210 33998 16213 34042
rect 16163 33995 16213 33998
rect 14913 33987 14971 33990
rect 14913 33935 14916 33987
rect 14968 33935 14971 33987
rect 14913 33932 14971 33935
rect 16163 33978 16213 33981
rect 16163 33934 16166 33978
rect 16210 33934 16213 33978
rect 16163 33931 16213 33934
rect 14897 33896 14929 33899
rect 14897 33838 14900 33896
rect 14926 33838 14929 33896
rect 14897 33835 14929 33838
rect 5090 33767 5141 33818
rect 3640 33760 5141 33767
rect 5167 33760 5170 33818
rect 14790 33760 14793 33818
rect 14819 33767 14870 33818
rect 16240 33767 16320 34125
rect 14819 33760 16320 33767
rect 3640 33725 5170 33760
rect 3000 33359 3003 33417
rect 3047 33359 3050 33417
rect 3000 33356 3050 33359
rect 3640 33367 3720 33725
rect 3747 33642 3797 33645
rect 3747 33598 3750 33642
rect 3794 33598 3797 33642
rect 3747 33595 3797 33598
rect 4989 33587 5047 33590
rect 3747 33578 3797 33581
rect 3747 33534 3750 33578
rect 3794 33534 3797 33578
rect 3747 33531 3797 33534
rect 4989 33535 4992 33587
rect 5044 33535 5047 33587
rect 4989 33532 5047 33535
rect 5031 33496 5063 33499
rect 5031 33438 5034 33496
rect 5060 33438 5063 33496
rect 5031 33435 5063 33438
rect 5090 33367 5170 33725
rect 14790 33725 16320 33760
rect 2936 31949 2939 32007
rect 2983 31949 2986 32007
rect 2936 31946 2986 31949
rect 3640 33325 5170 33367
rect 3640 32967 3720 33325
rect 3747 33242 3797 33245
rect 3747 33198 3750 33242
rect 3794 33198 3797 33242
rect 3747 33195 3797 33198
rect 4989 33187 5047 33190
rect 3747 33178 3797 33181
rect 3747 33134 3750 33178
rect 3794 33134 3797 33178
rect 3747 33131 3797 33134
rect 4989 33135 4992 33187
rect 5044 33135 5047 33187
rect 4989 33132 5047 33135
rect 5031 33096 5063 33099
rect 5031 33038 5034 33096
rect 5060 33038 5063 33096
rect 5031 33035 5063 33038
rect 5090 33018 5170 33325
rect 14790 33367 14870 33725
rect 16163 33642 16213 33645
rect 16163 33598 16166 33642
rect 16210 33598 16213 33642
rect 16163 33595 16213 33598
rect 14913 33587 14971 33590
rect 14913 33535 14916 33587
rect 14968 33535 14971 33587
rect 14913 33532 14971 33535
rect 16163 33578 16213 33581
rect 16163 33534 16166 33578
rect 16210 33534 16213 33578
rect 16163 33531 16213 33534
rect 14897 33496 14929 33499
rect 14897 33438 14900 33496
rect 14926 33438 14929 33496
rect 14897 33435 14929 33438
rect 16240 33367 16320 33725
rect 16846 33507 16896 38798
rect 16846 33449 16849 33507
rect 16893 33449 16896 33507
rect 16846 33446 16896 33449
rect 16910 38792 16960 38795
rect 16910 38734 16913 38792
rect 16957 38734 16960 38792
rect 14790 33325 16320 33367
rect 16910 33417 16960 38734
rect 16910 33359 16913 33417
rect 16957 33359 16960 33417
rect 16910 33356 16960 33359
rect 16974 38456 17024 38459
rect 16974 38398 16977 38456
rect 17021 38398 17024 38456
rect 14790 33018 14870 33325
rect 16163 33242 16213 33245
rect 16163 33198 16166 33242
rect 16210 33198 16213 33242
rect 16163 33195 16213 33198
rect 14913 33187 14971 33190
rect 14913 33135 14916 33187
rect 14968 33135 14971 33187
rect 14913 33132 14971 33135
rect 16163 33178 16213 33181
rect 16163 33134 16166 33178
rect 16210 33134 16213 33178
rect 16163 33131 16213 33134
rect 14897 33096 14929 33099
rect 14897 33038 14900 33096
rect 14926 33038 14929 33096
rect 14897 33035 14929 33038
rect 5090 32967 5141 33018
rect 3640 32960 5141 32967
rect 5167 32960 5170 33018
rect 14790 32960 14793 33018
rect 14819 32967 14870 33018
rect 16240 32967 16320 33325
rect 14819 32960 16320 32967
rect 3640 32925 5170 32960
rect 3640 32567 3720 32925
rect 3747 32842 3797 32845
rect 3747 32798 3750 32842
rect 3794 32798 3797 32842
rect 3747 32795 3797 32798
rect 4989 32787 5047 32790
rect 3747 32778 3797 32781
rect 3747 32734 3750 32778
rect 3794 32734 3797 32778
rect 3747 32731 3797 32734
rect 4989 32735 4992 32787
rect 5044 32735 5047 32787
rect 4989 32732 5047 32735
rect 5031 32696 5063 32699
rect 5031 32638 5034 32696
rect 5060 32638 5063 32696
rect 5031 32635 5063 32638
rect 5090 32567 5170 32925
rect 14790 32925 16320 32960
rect 3640 32525 5170 32567
rect 3640 32167 3720 32525
rect 3747 32442 3797 32445
rect 3747 32398 3750 32442
rect 3794 32398 3797 32442
rect 3747 32395 3797 32398
rect 4989 32387 5047 32390
rect 3747 32378 3797 32381
rect 3747 32334 3750 32378
rect 3794 32334 3797 32378
rect 3747 32331 3797 32334
rect 4989 32335 4992 32387
rect 5044 32335 5047 32387
rect 4989 32332 5047 32335
rect 5031 32296 5063 32299
rect 5031 32238 5034 32296
rect 5060 32238 5063 32296
rect 5031 32235 5063 32238
rect 5090 32218 5170 32525
rect 14790 32567 14870 32925
rect 16163 32842 16213 32845
rect 16163 32798 16166 32842
rect 16210 32798 16213 32842
rect 16163 32795 16213 32798
rect 14913 32787 14971 32790
rect 14913 32735 14916 32787
rect 14968 32735 14971 32787
rect 14913 32732 14971 32735
rect 16163 32778 16213 32781
rect 16163 32734 16166 32778
rect 16210 32734 16213 32778
rect 16163 32731 16213 32734
rect 14897 32696 14929 32699
rect 14897 32638 14900 32696
rect 14926 32638 14929 32696
rect 14897 32635 14929 32638
rect 16240 32567 16320 32925
rect 14790 32525 16320 32567
rect 14790 32218 14870 32525
rect 16163 32442 16213 32445
rect 16163 32398 16166 32442
rect 16210 32398 16213 32442
rect 16163 32395 16213 32398
rect 14913 32387 14971 32390
rect 14913 32335 14916 32387
rect 14968 32335 14971 32387
rect 14913 32332 14971 32335
rect 16163 32378 16213 32381
rect 16163 32334 16166 32378
rect 16210 32334 16213 32378
rect 16163 32331 16213 32334
rect 14897 32296 14929 32299
rect 14897 32238 14900 32296
rect 14926 32238 14929 32296
rect 14897 32235 14929 32238
rect 5090 32167 5141 32218
rect 3640 32160 5141 32167
rect 5167 32160 5170 32218
rect 14790 32160 14793 32218
rect 14819 32167 14870 32218
rect 16240 32167 16320 32525
rect 14819 32160 16320 32167
rect 3640 32125 5170 32160
rect 2872 31859 2875 31917
rect 2919 31859 2922 31917
rect 2872 31856 2922 31859
rect 2808 30449 2811 30507
rect 2855 30449 2858 30507
rect 2808 30446 2858 30449
rect 3640 31767 3720 32125
rect 3747 32042 3797 32045
rect 3747 31998 3750 32042
rect 3794 31998 3797 32042
rect 3747 31995 3797 31998
rect 4989 31987 5047 31990
rect 3747 31978 3797 31981
rect 3747 31934 3750 31978
rect 3794 31934 3797 31978
rect 3747 31931 3797 31934
rect 4989 31935 4992 31987
rect 5044 31935 5047 31987
rect 4989 31932 5047 31935
rect 5031 31896 5063 31899
rect 5031 31838 5034 31896
rect 5060 31838 5063 31896
rect 5031 31835 5063 31838
rect 5090 31767 5170 32125
rect 14790 32125 16320 32160
rect 3640 31725 5170 31767
rect 3640 31367 3720 31725
rect 3747 31642 3797 31645
rect 3747 31598 3750 31642
rect 3794 31598 3797 31642
rect 3747 31595 3797 31598
rect 4989 31587 5047 31590
rect 3747 31578 3797 31581
rect 3747 31534 3750 31578
rect 3794 31534 3797 31578
rect 3747 31531 3797 31534
rect 4989 31535 4992 31587
rect 5044 31535 5047 31587
rect 4989 31532 5047 31535
rect 5031 31496 5063 31499
rect 5031 31438 5034 31496
rect 5060 31438 5063 31496
rect 5031 31435 5063 31438
rect 5090 31418 5170 31725
rect 14790 31767 14870 32125
rect 16163 32042 16213 32045
rect 16163 31998 16166 32042
rect 16210 31998 16213 32042
rect 16163 31995 16213 31998
rect 14913 31987 14971 31990
rect 14913 31935 14916 31987
rect 14968 31935 14971 31987
rect 14913 31932 14971 31935
rect 16163 31978 16213 31981
rect 16163 31934 16166 31978
rect 16210 31934 16213 31978
rect 16163 31931 16213 31934
rect 14897 31896 14929 31899
rect 14897 31838 14900 31896
rect 14926 31838 14929 31896
rect 14897 31835 14929 31838
rect 16240 31767 16320 32125
rect 16974 32007 17024 38398
rect 16974 31949 16977 32007
rect 17021 31949 17024 32007
rect 16974 31946 17024 31949
rect 17038 38392 17088 38395
rect 17038 38334 17041 38392
rect 17085 38334 17088 38392
rect 17038 31917 17088 38334
rect 17038 31859 17041 31917
rect 17085 31859 17088 31917
rect 17038 31856 17088 31859
rect 17102 38155 17152 38158
rect 17102 38097 17105 38155
rect 17149 38097 17152 38155
rect 14790 31725 16320 31767
rect 14790 31418 14870 31725
rect 16163 31642 16213 31645
rect 16163 31598 16166 31642
rect 16210 31598 16213 31642
rect 16163 31595 16213 31598
rect 14913 31587 14971 31590
rect 14913 31535 14916 31587
rect 14968 31535 14971 31587
rect 14913 31532 14971 31535
rect 16163 31578 16213 31581
rect 16163 31534 16166 31578
rect 16210 31534 16213 31578
rect 16163 31531 16213 31534
rect 14897 31496 14929 31499
rect 14897 31438 14900 31496
rect 14926 31438 14929 31496
rect 14897 31435 14929 31438
rect 5090 31367 5141 31418
rect 3640 31360 5141 31367
rect 5167 31360 5170 31418
rect 14790 31360 14793 31418
rect 14819 31367 14870 31418
rect 16240 31367 16320 31725
rect 14819 31360 16320 31367
rect 3640 31325 5170 31360
rect 3640 30967 3720 31325
rect 3747 31242 3797 31245
rect 3747 31198 3750 31242
rect 3794 31198 3797 31242
rect 3747 31195 3797 31198
rect 4989 31187 5047 31190
rect 3747 31178 3797 31181
rect 3747 31134 3750 31178
rect 3794 31134 3797 31178
rect 3747 31131 3797 31134
rect 4989 31135 4992 31187
rect 5044 31135 5047 31187
rect 4989 31132 5047 31135
rect 5031 31096 5063 31099
rect 5031 31038 5034 31096
rect 5060 31038 5063 31096
rect 5031 31035 5063 31038
rect 5090 30967 5170 31325
rect 14790 31325 16320 31360
rect 3640 30925 5170 30967
rect 3640 30567 3720 30925
rect 3747 30842 3797 30845
rect 3747 30798 3750 30842
rect 3794 30798 3797 30842
rect 3747 30795 3797 30798
rect 4989 30787 5047 30790
rect 3747 30778 3797 30781
rect 3747 30734 3750 30778
rect 3794 30734 3797 30778
rect 3747 30731 3797 30734
rect 4989 30735 4992 30787
rect 5044 30735 5047 30787
rect 4989 30732 5047 30735
rect 5031 30696 5063 30699
rect 5031 30638 5034 30696
rect 5060 30638 5063 30696
rect 5031 30635 5063 30638
rect 5090 30618 5170 30925
rect 14790 30967 14870 31325
rect 16163 31242 16213 31245
rect 16163 31198 16166 31242
rect 16210 31198 16213 31242
rect 16163 31195 16213 31198
rect 14913 31187 14971 31190
rect 14913 31135 14916 31187
rect 14968 31135 14971 31187
rect 14913 31132 14971 31135
rect 16163 31178 16213 31181
rect 16163 31134 16166 31178
rect 16210 31134 16213 31178
rect 16163 31131 16213 31134
rect 14897 31096 14929 31099
rect 14897 31038 14900 31096
rect 14926 31038 14929 31096
rect 14897 31035 14929 31038
rect 16240 30967 16320 31325
rect 14790 30925 16320 30967
rect 14790 30618 14870 30925
rect 16163 30842 16213 30845
rect 16163 30798 16166 30842
rect 16210 30798 16213 30842
rect 16163 30795 16213 30798
rect 14913 30787 14971 30790
rect 14913 30735 14916 30787
rect 14968 30735 14971 30787
rect 14913 30732 14971 30735
rect 16163 30778 16213 30781
rect 16163 30734 16166 30778
rect 16210 30734 16213 30778
rect 16163 30731 16213 30734
rect 14897 30696 14929 30699
rect 14897 30638 14900 30696
rect 14926 30638 14929 30696
rect 14897 30635 14929 30638
rect 5090 30567 5141 30618
rect 3640 30560 5141 30567
rect 5167 30560 5170 30618
rect 14790 30560 14793 30618
rect 14819 30567 14870 30618
rect 16240 30567 16320 30925
rect 14819 30560 16320 30567
rect 3640 30525 5170 30560
rect 2744 30359 2747 30417
rect 2791 30359 2794 30417
rect 2744 30356 2794 30359
rect 2680 28949 2683 29007
rect 2727 28949 2730 29007
rect 2680 28946 2730 28949
rect 3640 30167 3720 30525
rect 3747 30442 3797 30445
rect 3747 30398 3750 30442
rect 3794 30398 3797 30442
rect 3747 30395 3797 30398
rect 4989 30387 5047 30390
rect 3747 30378 3797 30381
rect 3747 30334 3750 30378
rect 3794 30334 3797 30378
rect 3747 30331 3797 30334
rect 4989 30335 4992 30387
rect 5044 30335 5047 30387
rect 4989 30332 5047 30335
rect 5031 30296 5063 30299
rect 5031 30238 5034 30296
rect 5060 30238 5063 30296
rect 5031 30235 5063 30238
rect 5090 30167 5170 30525
rect 14790 30525 16320 30560
rect 3640 30125 5170 30167
rect 3640 29767 3720 30125
rect 3747 30042 3797 30045
rect 3747 29998 3750 30042
rect 3794 29998 3797 30042
rect 3747 29995 3797 29998
rect 4989 29987 5047 29990
rect 3747 29978 3797 29981
rect 3747 29934 3750 29978
rect 3794 29934 3797 29978
rect 3747 29931 3797 29934
rect 4989 29935 4992 29987
rect 5044 29935 5047 29987
rect 4989 29932 5047 29935
rect 5031 29896 5063 29899
rect 5031 29838 5034 29896
rect 5060 29838 5063 29896
rect 5031 29835 5063 29838
rect 5090 29818 5170 30125
rect 14790 30167 14870 30525
rect 16163 30442 16213 30445
rect 16163 30398 16166 30442
rect 16210 30398 16213 30442
rect 16163 30395 16213 30398
rect 14913 30387 14971 30390
rect 14913 30335 14916 30387
rect 14968 30335 14971 30387
rect 14913 30332 14971 30335
rect 16163 30378 16213 30381
rect 16163 30334 16166 30378
rect 16210 30334 16213 30378
rect 16163 30331 16213 30334
rect 14897 30296 14929 30299
rect 14897 30238 14900 30296
rect 14926 30238 14929 30296
rect 14897 30235 14929 30238
rect 16240 30167 16320 30525
rect 17102 30507 17152 38097
rect 17102 30449 17105 30507
rect 17149 30449 17152 30507
rect 17102 30446 17152 30449
rect 17166 38091 17216 38094
rect 17166 38033 17169 38091
rect 17213 38033 17216 38091
rect 17166 30417 17216 38033
rect 17166 30359 17169 30417
rect 17213 30359 17216 30417
rect 17166 30356 17216 30359
rect 17230 37656 17280 37659
rect 17230 37598 17233 37656
rect 17277 37598 17280 37656
rect 14790 30125 16320 30167
rect 14790 29818 14870 30125
rect 16163 30042 16213 30045
rect 16163 29998 16166 30042
rect 16210 29998 16213 30042
rect 16163 29995 16213 29998
rect 14913 29987 14971 29990
rect 14913 29935 14916 29987
rect 14968 29935 14971 29987
rect 14913 29932 14971 29935
rect 16163 29978 16213 29981
rect 16163 29934 16166 29978
rect 16210 29934 16213 29978
rect 16163 29931 16213 29934
rect 14897 29896 14929 29899
rect 14897 29838 14900 29896
rect 14926 29838 14929 29896
rect 14897 29835 14929 29838
rect 5090 29767 5141 29818
rect 3640 29760 5141 29767
rect 5167 29760 5170 29818
rect 14790 29760 14793 29818
rect 14819 29767 14870 29818
rect 16240 29767 16320 30125
rect 14819 29760 16320 29767
rect 3640 29725 5170 29760
rect 3640 29367 3720 29725
rect 3747 29642 3797 29645
rect 3747 29598 3750 29642
rect 3794 29598 3797 29642
rect 3747 29595 3797 29598
rect 4989 29587 5047 29590
rect 3747 29578 3797 29581
rect 3747 29534 3750 29578
rect 3794 29534 3797 29578
rect 3747 29531 3797 29534
rect 4989 29535 4992 29587
rect 5044 29535 5047 29587
rect 4989 29532 5047 29535
rect 5031 29496 5063 29499
rect 5031 29438 5034 29496
rect 5060 29438 5063 29496
rect 5031 29435 5063 29438
rect 5090 29367 5170 29725
rect 14790 29725 16320 29760
rect 3640 29325 5170 29367
rect 14790 29367 14870 29725
rect 16163 29642 16213 29645
rect 16163 29598 16166 29642
rect 16210 29598 16213 29642
rect 16163 29595 16213 29598
rect 14913 29587 14971 29590
rect 14913 29535 14916 29587
rect 14968 29535 14971 29587
rect 14913 29532 14971 29535
rect 16163 29578 16213 29581
rect 16163 29534 16166 29578
rect 16210 29534 16213 29578
rect 16163 29531 16213 29534
rect 14897 29496 14929 29499
rect 14897 29438 14900 29496
rect 14926 29438 14929 29496
rect 14897 29435 14929 29438
rect 16240 29367 16320 29725
rect 3640 28983 3720 29325
rect 3747 29242 3797 29245
rect 3747 29198 3750 29242
rect 3794 29198 3797 29242
rect 3747 29195 3797 29198
rect 4989 29187 5047 29190
rect 3747 29178 3797 29181
rect 3747 29134 3750 29178
rect 3794 29134 3797 29178
rect 3747 29131 3797 29134
rect 4989 29135 4992 29187
rect 5044 29135 5047 29187
rect 4989 29132 5047 29135
rect 5031 29096 5063 29099
rect 5031 29038 5034 29096
rect 5060 29038 5063 29096
rect 5031 29035 5063 29038
rect 5090 29000 5170 29325
rect 5210 29096 5290 29352
rect 5210 29038 5213 29096
rect 5239 29038 5290 29096
rect 5210 29035 5290 29038
rect 14670 29096 14750 29353
rect 14670 29038 14721 29096
rect 14747 29038 14750 29096
rect 14670 29035 14750 29038
rect 14790 29325 16320 29367
rect 14790 29000 14870 29325
rect 16163 29242 16213 29245
rect 16163 29198 16166 29242
rect 16210 29198 16213 29242
rect 16163 29195 16213 29198
rect 14913 29187 14971 29190
rect 14913 29135 14916 29187
rect 14968 29135 14971 29187
rect 14913 29132 14971 29135
rect 16163 29178 16213 29181
rect 16163 29134 16166 29178
rect 16210 29134 16213 29178
rect 16163 29131 16213 29134
rect 14897 29096 14929 29099
rect 14897 29038 14900 29096
rect 14926 29038 14929 29096
rect 14897 29035 14929 29038
rect 5090 28997 5820 29000
rect 5090 28983 5175 28997
rect 2616 28859 2619 28917
rect 2663 28859 2666 28917
rect 3640 28908 5175 28983
rect 5815 28908 5820 28997
rect 3640 28903 5820 28908
rect 14140 28997 14870 29000
rect 14140 28908 14145 28997
rect 14785 28983 14870 28997
rect 16240 28983 16320 29325
rect 14785 28908 16320 28983
rect 17230 29007 17280 37598
rect 17230 28949 17233 29007
rect 17277 28949 17280 29007
rect 17230 28946 17280 28949
rect 17294 37592 17344 37595
rect 17294 37534 17297 37592
rect 17341 37534 17344 37592
rect 14140 28903 16320 28908
rect 17294 28917 17344 37534
rect 2616 28856 2666 28859
rect 17294 28859 17297 28917
rect 17341 28859 17344 28917
rect 17294 28856 17344 28859
rect 17358 37256 17408 37259
rect 17358 37198 17361 37256
rect 17405 37198 17408 37256
rect 2552 27449 2555 27507
rect 2599 27449 2602 27507
rect 2552 27446 2602 27449
rect 17358 27507 17408 37198
rect 17358 27449 17361 27507
rect 17405 27449 17408 27507
rect 17358 27446 17408 27449
rect 17422 37192 17472 37195
rect 17422 37134 17425 37192
rect 17469 37134 17472 37192
rect 2488 27359 2491 27417
rect 2535 27359 2538 27417
rect 2488 27356 2538 27359
rect 17422 27417 17472 37134
rect 17422 27359 17425 27417
rect 17469 27359 17472 27417
rect 17422 27356 17472 27359
rect 17486 36856 17536 36859
rect 17486 36798 17489 36856
rect 17533 36798 17536 36856
rect 2424 25949 2427 26007
rect 2471 25949 2474 26007
rect 2424 25946 2474 25949
rect 17486 26007 17536 36798
rect 17486 25949 17489 26007
rect 17533 25949 17536 26007
rect 17486 25946 17536 25949
rect 17550 36792 17600 36795
rect 17550 36734 17553 36792
rect 17597 36734 17600 36792
rect 2360 25859 2363 25917
rect 2407 25859 2410 25917
rect 2360 25856 2410 25859
rect 17550 25917 17600 36734
rect 17550 25859 17553 25917
rect 17597 25859 17600 25917
rect 17550 25856 17600 25859
rect 17614 36655 17664 36658
rect 17614 36597 17617 36655
rect 17661 36597 17664 36655
rect 2296 24449 2299 24507
rect 2343 24449 2346 24507
rect 2296 24446 2346 24449
rect 17614 24507 17664 36597
rect 17614 24449 17617 24507
rect 17661 24449 17664 24507
rect 17614 24446 17664 24449
rect 17678 36591 17728 36594
rect 17678 36533 17681 36591
rect 17725 36533 17728 36591
rect 2232 24359 2235 24417
rect 2279 24359 2282 24417
rect 2232 24356 2282 24359
rect 17678 24417 17728 36533
rect 17678 24359 17681 24417
rect 17725 24359 17728 24417
rect 17678 24356 17728 24359
rect 17742 36056 17792 36059
rect 17742 35998 17745 36056
rect 17789 35998 17792 36056
rect 2168 22949 2171 23007
rect 2215 22949 2218 23007
rect 2168 22946 2218 22949
rect 17742 23007 17792 35998
rect 17742 22949 17745 23007
rect 17789 22949 17792 23007
rect 17742 22946 17792 22949
rect 17806 35992 17856 35995
rect 17806 35934 17809 35992
rect 17853 35934 17856 35992
rect 2104 22859 2107 22917
rect 2151 22859 2154 22917
rect 2104 22856 2154 22859
rect 17806 22917 17856 35934
rect 17806 22859 17809 22917
rect 17853 22859 17856 22917
rect 17806 22856 17856 22859
rect 17870 35656 17920 35659
rect 17870 35598 17873 35656
rect 17917 35598 17920 35656
rect 2040 21449 2043 21507
rect 2087 21449 2090 21507
rect 2040 21446 2090 21449
rect 17870 21507 17920 35598
rect 17870 21449 17873 21507
rect 17917 21449 17920 21507
rect 17870 21446 17920 21449
rect 17934 35592 17984 35595
rect 17934 35534 17937 35592
rect 17981 35534 17984 35592
rect 1976 21359 1979 21417
rect 2023 21359 2026 21417
rect 1976 21356 2026 21359
rect 17934 21417 17984 35534
rect 17934 21359 17937 21417
rect 17981 21359 17984 21417
rect 17934 21356 17984 21359
rect 17998 35256 18048 35259
rect 17998 35198 18001 35256
rect 18045 35198 18048 35256
rect 1912 19949 1915 20007
rect 1959 19949 1962 20007
rect 1912 19946 1962 19949
rect 17998 20007 18048 35198
rect 17998 19949 18001 20007
rect 18045 19949 18048 20007
rect 17998 19946 18048 19949
rect 18062 35192 18112 35195
rect 18062 35134 18065 35192
rect 18109 35134 18112 35192
rect 1848 19859 1851 19917
rect 1895 19859 1898 19917
rect 1848 19856 1898 19859
rect 18062 19917 18112 35134
rect 18062 19859 18065 19917
rect 18109 19859 18112 19917
rect 18062 19856 18112 19859
rect 18126 34853 18176 34856
rect 18126 34795 18129 34853
rect 18173 34795 18176 34853
rect 1784 18449 1787 18507
rect 1831 18449 1834 18507
rect 1784 18446 1834 18449
rect 18126 18507 18176 34795
rect 18126 18449 18129 18507
rect 18173 18449 18176 18507
rect 18126 18446 18176 18449
rect 18190 34789 18240 34792
rect 18190 34731 18193 34789
rect 18237 34731 18240 34789
rect 1720 18359 1723 18417
rect 1767 18359 1770 18417
rect 1720 18356 1770 18359
rect 18190 18417 18240 34731
rect 18190 18359 18193 18417
rect 18237 18359 18240 18417
rect 18190 18356 18240 18359
rect 18254 34456 18304 34459
rect 18254 34398 18257 34456
rect 18301 34398 18304 34456
rect 1656 16949 1659 17007
rect 1703 16949 1706 17007
rect 1656 16946 1706 16949
rect 18254 17007 18304 34398
rect 18254 16949 18257 17007
rect 18301 16949 18304 17007
rect 18254 16946 18304 16949
rect 18318 34392 18368 34395
rect 18318 34334 18321 34392
rect 18365 34334 18368 34392
rect 1592 16859 1595 16917
rect 1639 16859 1642 16917
rect 1592 16856 1642 16859
rect 18318 16917 18368 34334
rect 18318 16859 18321 16917
rect 18365 16859 18368 16917
rect 18318 16856 18368 16859
rect 18382 34056 18432 34059
rect 18382 33998 18385 34056
rect 18429 33998 18432 34056
rect 1528 15449 1531 15507
rect 1575 15449 1578 15507
rect 1528 15446 1578 15449
rect 18382 15507 18432 33998
rect 18382 15449 18385 15507
rect 18429 15449 18432 15507
rect 18382 15446 18432 15449
rect 18446 33992 18496 33995
rect 18446 33934 18449 33992
rect 18493 33934 18496 33992
rect 1464 15359 1467 15417
rect 1511 15359 1514 15417
rect 1464 15356 1514 15359
rect 18446 15417 18496 33934
rect 18446 15359 18449 15417
rect 18493 15359 18496 15417
rect 18446 15356 18496 15359
rect 18510 33656 18560 33659
rect 18510 33598 18513 33656
rect 18557 33598 18560 33656
rect 1400 13949 1403 14007
rect 1447 13949 1450 14007
rect 1400 13946 1450 13949
rect 18510 14007 18560 33598
rect 18510 13949 18513 14007
rect 18557 13949 18560 14007
rect 18510 13946 18560 13949
rect 18574 33592 18624 33595
rect 18574 33534 18577 33592
rect 18621 33534 18624 33592
rect 1336 13859 1339 13917
rect 1383 13859 1386 13917
rect 1336 13856 1386 13859
rect 18574 13917 18624 33534
rect 18574 13859 18577 13917
rect 18621 13859 18624 13917
rect 18574 13856 18624 13859
rect 18638 33256 18688 33259
rect 18638 33198 18641 33256
rect 18685 33198 18688 33256
rect 1272 12449 1275 12507
rect 1319 12449 1322 12507
rect 1272 12446 1322 12449
rect 18638 12507 18688 33198
rect 18638 12449 18641 12507
rect 18685 12449 18688 12507
rect 18638 12446 18688 12449
rect 18702 33192 18752 33195
rect 18702 33134 18705 33192
rect 18749 33134 18752 33192
rect 1208 12359 1211 12417
rect 1255 12359 1258 12417
rect 1208 12356 1258 12359
rect 18702 12417 18752 33134
rect 18702 12359 18705 12417
rect 18749 12359 18752 12417
rect 18702 12356 18752 12359
rect 18766 32856 18816 32859
rect 18766 32798 18769 32856
rect 18813 32798 18816 32856
rect 1144 10949 1147 11007
rect 1191 10949 1194 11007
rect 1144 10946 1194 10949
rect 18766 11007 18816 32798
rect 18766 10949 18769 11007
rect 18813 10949 18816 11007
rect 18766 10946 18816 10949
rect 18830 32792 18880 32795
rect 18830 32734 18833 32792
rect 18877 32734 18880 32792
rect 1080 10859 1083 10917
rect 1127 10859 1130 10917
rect 1080 10856 1130 10859
rect 18830 10917 18880 32734
rect 18830 10859 18833 10917
rect 18877 10859 18880 10917
rect 18830 10856 18880 10859
rect 18894 32456 18944 32459
rect 18894 32398 18897 32456
rect 18941 32398 18944 32456
rect 1016 9449 1019 9507
rect 1063 9449 1066 9507
rect 1016 9446 1066 9449
rect 18894 9507 18944 32398
rect 18894 9449 18897 9507
rect 18941 9449 18944 9507
rect 18894 9446 18944 9449
rect 18958 32392 19008 32395
rect 18958 32334 18961 32392
rect 19005 32334 19008 32392
rect 952 9359 955 9417
rect 999 9359 1002 9417
rect 952 9356 1002 9359
rect 18958 9417 19008 32334
rect 18958 9359 18961 9417
rect 19005 9359 19008 9417
rect 18958 9356 19008 9359
rect 19022 32149 19072 32152
rect 19022 32091 19025 32149
rect 19069 32091 19072 32149
rect 888 7949 891 8007
rect 935 7949 938 8007
rect 888 7946 938 7949
rect 19022 8007 19072 32091
rect 19022 7949 19025 8007
rect 19069 7949 19072 8007
rect 19022 7946 19072 7949
rect 19086 32085 19136 32088
rect 19086 32027 19089 32085
rect 19133 32027 19136 32085
rect 824 7859 827 7917
rect 871 7859 874 7917
rect 824 7856 874 7859
rect 19086 7917 19136 32027
rect 19086 7859 19089 7917
rect 19133 7859 19136 7917
rect 19086 7856 19136 7859
rect 19150 31656 19200 31659
rect 19150 31598 19153 31656
rect 19197 31598 19200 31656
rect 760 6449 763 6507
rect 807 6449 810 6507
rect 760 6446 810 6449
rect 19150 6507 19200 31598
rect 19150 6449 19153 6507
rect 19197 6449 19200 6507
rect 19150 6446 19200 6449
rect 19214 31592 19264 31595
rect 19214 31534 19217 31592
rect 19261 31534 19264 31592
rect 696 6359 699 6417
rect 743 6359 746 6417
rect 696 6356 746 6359
rect 19214 6417 19264 31534
rect 19214 6359 19217 6417
rect 19261 6359 19264 6417
rect 19214 6356 19264 6359
rect 19278 31256 19328 31259
rect 19278 31198 19281 31256
rect 19325 31198 19328 31256
rect 12868 6201 12968 6204
rect 12868 6107 12871 6201
rect 12965 6107 12968 6201
rect 12868 5577 12968 6107
rect 12868 5483 12871 5577
rect 12965 5483 12968 5577
rect 12868 5480 12968 5483
rect 13006 6033 13106 6036
rect 13006 5939 13009 6033
rect 13103 5939 13106 6033
rect 13006 5577 13106 5939
rect 13006 5483 13009 5577
rect 13103 5483 13106 5577
rect 13006 5480 13106 5483
rect 13144 5865 13244 5868
rect 13144 5771 13147 5865
rect 13241 5771 13244 5865
rect 13144 5577 13244 5771
rect 13144 5483 13147 5577
rect 13241 5483 13244 5577
rect 13144 5480 13244 5483
rect 13282 5697 13382 5700
rect 13282 5603 13285 5697
rect 13379 5603 13382 5697
rect 13282 5577 13382 5603
rect 13282 5483 13285 5577
rect 13379 5483 13382 5577
rect 13282 5480 13382 5483
rect 632 4949 635 5007
rect 679 4949 682 5007
rect 632 4946 682 4949
rect 19278 5007 19328 31198
rect 19278 4949 19281 5007
rect 19325 4949 19328 5007
rect 19278 4946 19328 4949
rect 19342 31192 19392 31195
rect 19342 31134 19345 31192
rect 19389 31134 19392 31192
rect 568 4859 571 4917
rect 615 4859 618 4917
rect 568 4856 618 4859
rect 19342 4917 19392 31134
rect 19342 4859 19345 4917
rect 19389 4859 19392 4917
rect 19342 4856 19392 4859
rect 19406 30856 19456 30859
rect 19406 30798 19409 30856
rect 19453 30798 19456 30856
rect 504 3449 507 3507
rect 551 3449 554 3507
rect 504 3446 554 3449
rect 19406 3507 19456 30798
rect 19406 3449 19409 3507
rect 19453 3449 19456 3507
rect 19406 3446 19456 3449
rect 19470 30792 19520 30795
rect 19470 30734 19473 30792
rect 19517 30734 19520 30792
rect 440 3359 443 3417
rect 487 3359 490 3417
rect 440 3356 490 3359
rect 19470 3417 19520 30734
rect 19470 3359 19473 3417
rect 19517 3359 19520 3417
rect 19470 3356 19520 3359
rect 19534 30655 19584 30658
rect 19534 30597 19537 30655
rect 19581 30597 19584 30655
rect 376 1949 379 2007
rect 423 1949 426 2007
rect 376 1946 426 1949
rect 5903 2541 6000 2630
rect 5903 1980 5983 2541
rect 6083 2049 6400 2100
rect 6083 2023 6086 2049
rect 6138 2023 6400 2049
rect 6083 2020 6400 2023
rect 19534 2007 19584 30597
rect 5903 1977 12520 1980
rect 5903 1951 6814 1977
rect 6866 1951 7614 1977
rect 7666 1951 8414 1977
rect 8466 1951 9214 1977
rect 9266 1951 10014 1977
rect 10066 1951 10814 1977
rect 10866 1951 11614 1977
rect 11666 1951 12443 1977
rect 312 1859 315 1917
rect 359 1859 362 1917
rect 5903 1903 12443 1951
rect 12517 1903 12520 1977
rect 19534 1949 19537 2007
rect 19581 1949 19584 2007
rect 19534 1946 19584 1949
rect 19598 30591 19648 30594
rect 19598 30533 19601 30591
rect 19645 30533 19648 30591
rect 5903 1900 12520 1903
rect 19598 1917 19648 30533
rect 312 1856 362 1859
rect 6083 1870 6141 1873
rect 6083 1844 6086 1870
rect 6138 1844 6141 1870
rect 6373 1867 6396 1900
rect 6483 1870 6541 1873
rect 6083 1841 6141 1844
rect 6483 1844 6486 1870
rect 6538 1844 6541 1870
rect 6773 1867 6796 1900
rect 6883 1870 6941 1873
rect 6483 1841 6541 1844
rect 6883 1844 6886 1870
rect 6938 1844 6941 1870
rect 7173 1867 7196 1900
rect 7283 1870 7341 1873
rect 6883 1841 6941 1844
rect 7283 1844 7286 1870
rect 7338 1844 7341 1870
rect 7573 1867 7596 1900
rect 7683 1870 7741 1873
rect 7283 1841 7341 1844
rect 7683 1844 7686 1870
rect 7738 1844 7741 1870
rect 7973 1867 7996 1900
rect 8083 1870 8141 1873
rect 7683 1841 7741 1844
rect 8083 1844 8086 1870
rect 8138 1844 8141 1870
rect 8373 1867 8396 1900
rect 8483 1870 8541 1873
rect 8083 1841 8141 1844
rect 8483 1844 8486 1870
rect 8538 1844 8541 1870
rect 8773 1867 8796 1900
rect 8883 1870 8941 1873
rect 8483 1841 8541 1844
rect 8883 1844 8886 1870
rect 8938 1844 8941 1870
rect 9173 1867 9196 1900
rect 9283 1870 9341 1873
rect 8883 1841 8941 1844
rect 9283 1844 9286 1870
rect 9338 1844 9341 1870
rect 9573 1867 9596 1900
rect 9683 1870 9741 1873
rect 9283 1841 9341 1844
rect 9683 1844 9686 1870
rect 9738 1844 9741 1870
rect 9973 1867 9996 1900
rect 10083 1870 10141 1873
rect 9683 1841 9741 1844
rect 10083 1844 10086 1870
rect 10138 1844 10141 1870
rect 10373 1867 10396 1900
rect 10483 1870 10541 1873
rect 10083 1841 10141 1844
rect 10483 1844 10486 1870
rect 10538 1844 10541 1870
rect 10773 1867 10796 1900
rect 10883 1870 10941 1873
rect 10483 1841 10541 1844
rect 10883 1844 10886 1870
rect 10938 1844 10941 1870
rect 11173 1867 11196 1900
rect 11283 1870 11341 1873
rect 10883 1841 10941 1844
rect 11283 1844 11286 1870
rect 11338 1844 11341 1870
rect 11573 1867 11596 1900
rect 11683 1870 11741 1873
rect 11283 1841 11341 1844
rect 11683 1844 11686 1870
rect 11738 1844 11741 1870
rect 11973 1867 11996 1900
rect 12083 1870 12141 1873
rect 11683 1841 11741 1844
rect 12083 1844 12086 1870
rect 12138 1844 12141 1870
rect 12373 1867 12396 1900
rect 19598 1859 19601 1917
rect 19645 1859 19648 1917
rect 19598 1856 19648 1859
rect 19662 30056 19712 30059
rect 19662 29998 19665 30056
rect 19709 29998 19712 30056
rect 12083 1841 12141 1844
rect 248 449 251 507
rect 295 449 298 507
rect 248 446 298 449
rect 184 359 187 417
rect 231 359 234 417
rect 184 356 234 359
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -220 -5 -140 0
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect -220 -80 -140 -75
rect -18268 -984 -18236 -981
rect -18268 -1010 -18265 -984
rect -18239 -1010 -18236 -984
rect -18268 -1018 -18236 -1010
rect -18206 -1018 -18156 -80
rect -16268 -892 -16236 -889
rect -16268 -918 -16265 -892
rect -16239 -918 -16236 -892
rect -18014 -938 -17982 -935
rect -18014 -964 -18011 -938
rect -17985 -964 -17982 -938
rect -18014 -1018 -17982 -964
rect -16268 -1018 -16236 -918
rect -16206 -1018 -16156 -80
rect -14268 -800 -14236 -797
rect -14268 -826 -14265 -800
rect -14239 -826 -14236 -800
rect -16014 -846 -15982 -843
rect -16014 -872 -16011 -846
rect -15985 -872 -15982 -846
rect -16014 -1018 -15982 -872
rect -14268 -1018 -14236 -826
rect -14206 -1018 -14156 -80
rect -12268 -708 -12236 -705
rect -12268 -734 -12265 -708
rect -12239 -734 -12236 -708
rect -14014 -754 -13982 -751
rect -14014 -780 -14011 -754
rect -13985 -780 -13982 -754
rect -14014 -1018 -13982 -780
rect -12268 -1018 -12236 -734
rect -12206 -1018 -12156 -80
rect -10268 -616 -10236 -613
rect -10268 -642 -10265 -616
rect -10239 -642 -10236 -616
rect -12014 -662 -11982 -659
rect -12014 -688 -12011 -662
rect -11985 -688 -11982 -662
rect -12014 -1018 -11982 -688
rect -10268 -1018 -10236 -642
rect -10206 -1018 -10156 -80
rect -8268 -524 -8236 -521
rect -8268 -550 -8265 -524
rect -8239 -550 -8236 -524
rect -10014 -570 -9982 -567
rect -10014 -596 -10011 -570
rect -9985 -596 -9982 -570
rect -10014 -1018 -9982 -596
rect -8268 -1018 -8236 -550
rect -8206 -1018 -8156 -80
rect -6268 -432 -6236 -429
rect -6268 -458 -6265 -432
rect -6239 -458 -6236 -432
rect -8014 -478 -7982 -475
rect -8014 -504 -8011 -478
rect -7985 -504 -7982 -478
rect -8014 -1018 -7982 -504
rect -6268 -1018 -6236 -458
rect -6206 -1018 -6156 -80
rect -4268 -340 -4236 -337
rect -4268 -366 -4265 -340
rect -4239 -366 -4236 -340
rect -6014 -386 -5982 -383
rect -6014 -412 -6011 -386
rect -5985 -412 -5982 -386
rect -6014 -1018 -5982 -412
rect -4268 -1018 -4236 -366
rect -4206 -1018 -4156 -80
rect -2268 -248 -2236 -245
rect -2268 -274 -2265 -248
rect -2239 -274 -2236 -248
rect -4014 -294 -3982 -291
rect -4014 -320 -4011 -294
rect -3985 -320 -3982 -294
rect -4014 -1018 -3982 -320
rect -2268 -1018 -2236 -274
rect -2206 -1018 -2156 -80
rect -268 -156 -236 -153
rect -268 -182 -265 -156
rect -239 -182 -236 -156
rect -2014 -202 -1982 -199
rect -2014 -228 -2011 -202
rect -1985 -228 -1982 -202
rect -2014 -1018 -1982 -228
rect -268 -1018 -236 -182
rect -206 -1018 -156 -80
rect -14 -110 18 -107
rect -14 -136 -11 -110
rect 15 -136 18 -110
rect -14 -1018 18 -136
rect 8593 -984 8625 557
rect 8647 -938 8679 557
rect 8993 -892 9025 557
rect 9047 -846 9079 557
rect 9393 -800 9425 557
rect 9447 -754 9479 557
rect 9793 -708 9825 557
rect 9847 -662 9879 557
rect 10193 -616 10225 557
rect 10247 -570 10279 557
rect 10593 -524 10625 557
rect 10647 -478 10679 557
rect 10993 -432 11025 557
rect 11047 -386 11079 557
rect 11393 -340 11425 557
rect 11447 -294 11479 557
rect 11793 -248 11825 557
rect 11847 -202 11879 557
rect 12193 -156 12225 557
rect 12247 -110 12279 557
rect 19662 507 19712 29998
rect 19662 449 19665 507
rect 19709 449 19712 507
rect 19662 446 19712 449
rect 19726 29992 19776 29995
rect 19726 29934 19729 29992
rect 19773 29934 19776 29992
rect 19726 417 19776 29934
rect 19726 359 19729 417
rect 19773 359 19776 417
rect 19726 356 19776 359
rect 20100 -5 20180 0
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
rect 12247 -136 12250 -110
rect 12276 -136 12279 -110
rect 12247 -139 12279 -136
rect 19941 -110 19973 -107
rect 19941 -136 19944 -110
rect 19970 -136 19973 -110
rect 12193 -182 12196 -156
rect 12222 -182 12225 -156
rect 12193 -185 12225 -182
rect 11847 -228 11850 -202
rect 11876 -228 11879 -202
rect 11847 -231 11879 -228
rect 11793 -274 11796 -248
rect 11822 -274 11825 -248
rect 11793 -277 11825 -274
rect 11447 -320 11450 -294
rect 11476 -320 11479 -294
rect 11447 -323 11479 -320
rect 11393 -366 11396 -340
rect 11422 -366 11425 -340
rect 11393 -369 11425 -366
rect 11047 -412 11050 -386
rect 11076 -412 11079 -386
rect 11047 -415 11079 -412
rect 10993 -458 10996 -432
rect 11022 -458 11025 -432
rect 10993 -461 11025 -458
rect 10647 -504 10650 -478
rect 10676 -504 10679 -478
rect 10647 -507 10679 -504
rect 10593 -550 10596 -524
rect 10622 -550 10625 -524
rect 10593 -553 10625 -550
rect 10247 -596 10250 -570
rect 10276 -596 10279 -570
rect 10247 -599 10279 -596
rect 10193 -642 10196 -616
rect 10222 -642 10225 -616
rect 10193 -645 10225 -642
rect 9847 -688 9850 -662
rect 9876 -688 9879 -662
rect 9847 -691 9879 -688
rect 9793 -734 9796 -708
rect 9822 -734 9825 -708
rect 9793 -737 9825 -734
rect 9447 -780 9450 -754
rect 9476 -780 9479 -754
rect 9447 -783 9479 -780
rect 9393 -826 9396 -800
rect 9422 -826 9425 -800
rect 9393 -829 9425 -826
rect 9047 -872 9050 -846
rect 9076 -872 9079 -846
rect 9047 -875 9079 -872
rect 8993 -918 8996 -892
rect 9022 -918 9025 -892
rect 8993 -921 9025 -918
rect 8647 -964 8650 -938
rect 8676 -964 8679 -938
rect 8647 -967 8679 -964
rect 8593 -1010 8596 -984
rect 8622 -1010 8625 -984
rect 8593 -1013 8625 -1010
rect 19941 -1018 19973 -136
rect 20115 -1018 20165 -80
rect 20195 -156 20227 -153
rect 20195 -182 20198 -156
rect 20224 -182 20227 -156
rect 20195 -1018 20227 -182
rect 21941 -202 21973 -199
rect 21941 -228 21944 -202
rect 21970 -228 21973 -202
rect 21941 -1018 21973 -228
rect 22115 -1018 22165 -80
rect 22195 -248 22227 -245
rect 22195 -274 22198 -248
rect 22224 -274 22227 -248
rect 22195 -1018 22227 -274
rect 23941 -294 23973 -291
rect 23941 -320 23944 -294
rect 23970 -320 23973 -294
rect 23941 -1018 23973 -320
rect 24115 -1018 24165 -80
rect 24195 -340 24227 -337
rect 24195 -366 24198 -340
rect 24224 -366 24227 -340
rect 24195 -1018 24227 -366
rect 25941 -386 25973 -383
rect 25941 -412 25944 -386
rect 25970 -412 25973 -386
rect 25941 -1018 25973 -412
rect 26115 -1018 26165 -80
rect 26195 -432 26227 -429
rect 26195 -458 26198 -432
rect 26224 -458 26227 -432
rect 26195 -1018 26227 -458
rect 27941 -478 27973 -475
rect 27941 -504 27944 -478
rect 27970 -504 27973 -478
rect 27941 -1018 27973 -504
rect 28115 -1018 28165 -80
rect 28195 -524 28227 -521
rect 28195 -550 28198 -524
rect 28224 -550 28227 -524
rect 28195 -1018 28227 -550
rect 29941 -570 29973 -567
rect 29941 -596 29944 -570
rect 29970 -596 29973 -570
rect 29941 -1018 29973 -596
rect 30115 -1018 30165 -80
rect 30195 -616 30227 -613
rect 30195 -642 30198 -616
rect 30224 -642 30227 -616
rect 30195 -1018 30227 -642
rect 31941 -662 31973 -659
rect 31941 -688 31944 -662
rect 31970 -688 31973 -662
rect 31941 -1018 31973 -688
rect 32115 -1018 32165 -80
rect 32195 -708 32227 -705
rect 32195 -734 32198 -708
rect 32224 -734 32227 -708
rect 32195 -1018 32227 -734
rect 33941 -754 33973 -751
rect 33941 -780 33944 -754
rect 33970 -780 33973 -754
rect 33941 -1018 33973 -780
rect 34115 -1018 34165 -80
rect 34195 -800 34227 -797
rect 34195 -826 34198 -800
rect 34224 -826 34227 -800
rect 34195 -1018 34227 -826
rect 35941 -846 35973 -843
rect 35941 -872 35944 -846
rect 35970 -872 35973 -846
rect 35941 -1018 35973 -872
rect 36115 -1018 36165 -80
rect 36195 -892 36227 -889
rect 36195 -918 36198 -892
rect 36224 -918 36227 -892
rect 36195 -1018 36227 -918
rect 37941 -938 37973 -935
rect 37941 -964 37944 -938
rect 37970 -964 37973 -938
rect 37941 -1018 37973 -964
rect 38115 -1018 38165 -80
rect 38195 -984 38227 -981
rect 38195 -1010 38198 -984
rect 38224 -1010 38227 -984
rect 38195 -1018 38227 -1010
<< via1 >>
rect 3259 43963 3303 44021
rect 16657 43963 16701 44021
rect 3259 41584 3303 41642
rect 3323 43873 3367 43931
rect 16593 43873 16637 43931
rect 3323 41520 3367 41578
rect 3387 42463 3431 42521
rect 16529 42463 16573 42521
rect 3387 41184 3431 41242
rect 3451 42373 3495 42431
rect 16465 42373 16509 42431
rect 3451 41120 3495 41178
rect 5090 41793 5170 41871
rect 14790 41793 14870 41871
rect 3750 41598 3794 41642
rect 3750 41534 3794 41578
rect 4992 41535 5044 41587
rect 5034 41438 5060 41496
rect 5213 41438 5239 41496
rect 14721 41438 14747 41496
rect 3515 40963 3559 41021
rect 3750 41198 3794 41242
rect 3750 41134 3794 41178
rect 4992 41135 5044 41187
rect 5034 41038 5060 41096
rect 16166 41598 16210 41642
rect 14916 41535 14968 41587
rect 16166 41534 16210 41578
rect 14900 41438 14926 41496
rect 5213 41038 5239 41096
rect 14721 41038 14747 41096
rect 16166 41198 16210 41242
rect 14916 41135 14968 41187
rect 16166 41134 16210 41178
rect 14900 41038 14926 41096
rect 5141 40960 5167 41018
rect 5320 40960 5346 41018
rect 14614 40960 14640 41018
rect 14793 40960 14819 41018
rect 16657 41584 16701 41642
rect 16593 41520 16637 41578
rect 16529 41184 16573 41242
rect 16465 41120 16509 41178
rect 3515 40784 3559 40842
rect 3579 40873 3623 40931
rect 3579 40720 3623 40778
rect 3750 40798 3794 40842
rect 3750 40734 3794 40778
rect 4992 40735 5044 40787
rect 5034 40638 5060 40696
rect 16401 40963 16445 41021
rect 5213 40638 5239 40696
rect 14721 40638 14747 40696
rect 3579 40398 3623 40456
rect 3515 40334 3559 40392
rect 3451 39998 3495 40056
rect 3387 39934 3431 39992
rect 3323 39598 3367 39656
rect 3259 39534 3303 39592
rect 3195 39198 3239 39256
rect 3131 39134 3175 39192
rect 3067 38798 3111 38856
rect 3003 38734 3047 38792
rect 2939 38398 2983 38456
rect 2875 38334 2919 38392
rect 2811 38097 2855 38155
rect 2747 38033 2791 38091
rect 2683 37598 2727 37656
rect 2619 37534 2663 37592
rect 2555 37198 2599 37256
rect 2491 37134 2535 37192
rect 2427 36798 2471 36856
rect 2363 36734 2407 36792
rect 2299 36597 2343 36655
rect 2235 36533 2279 36591
rect 2171 35998 2215 36056
rect 2107 35934 2151 35992
rect 2043 35598 2087 35656
rect 1979 35534 2023 35592
rect 1915 35198 1959 35256
rect 1851 35134 1895 35192
rect 1787 34795 1831 34853
rect 1723 34731 1767 34789
rect 1659 34398 1703 34456
rect 1595 34334 1639 34392
rect 1531 33998 1575 34056
rect 1467 33934 1511 33992
rect 1403 33598 1447 33656
rect 1339 33534 1383 33592
rect 1275 33198 1319 33256
rect 1211 33134 1255 33192
rect 1147 32798 1191 32856
rect 1083 32734 1127 32792
rect 1019 32398 1063 32456
rect 955 32334 999 32392
rect 891 32091 935 32149
rect 827 32027 871 32085
rect 763 31598 807 31656
rect 699 31534 743 31592
rect 635 31198 679 31256
rect 571 31134 615 31192
rect 507 30798 551 30856
rect 443 30734 487 30792
rect 379 30597 423 30655
rect 315 30533 359 30591
rect 251 29998 295 30056
rect 187 29934 231 29992
rect 3579 39449 3623 39507
rect 3750 40398 3794 40442
rect 3750 40334 3794 40378
rect 4992 40335 5044 40387
rect 5034 40238 5060 40296
rect 16166 40798 16210 40842
rect 14916 40735 14968 40787
rect 16166 40734 16210 40778
rect 14900 40638 14926 40696
rect 16337 40873 16381 40931
rect 16401 40784 16445 40842
rect 16337 40720 16381 40778
rect 5213 40238 5239 40296
rect 14721 40238 14747 40296
rect 16166 40398 16210 40442
rect 14916 40335 14968 40387
rect 16166 40334 16210 40378
rect 14900 40238 14926 40296
rect 5141 40160 5167 40218
rect 5320 40160 5346 40218
rect 14614 40160 14640 40218
rect 14793 40160 14819 40218
rect 3750 39998 3794 40042
rect 3750 39934 3794 39978
rect 4992 39935 5044 39987
rect 5034 39838 5060 39896
rect 5213 39838 5239 39896
rect 14721 39838 14747 39896
rect 3515 39359 3559 39417
rect 3750 39598 3794 39642
rect 3750 39534 3794 39578
rect 4992 39535 5044 39587
rect 5034 39438 5060 39496
rect 16166 39998 16210 40042
rect 14916 39935 14968 39987
rect 16166 39934 16210 39978
rect 14900 39838 14926 39896
rect 5213 39438 5239 39496
rect 14721 39438 14747 39496
rect 16166 39598 16210 39642
rect 14916 39535 14968 39587
rect 16166 39534 16210 39578
rect 14900 39438 14926 39496
rect 5141 39360 5167 39418
rect 5320 39360 5346 39418
rect 14614 39360 14640 39418
rect 14793 39360 14819 39418
rect 16337 40398 16381 40456
rect 16337 39449 16381 39507
rect 16401 40334 16445 40392
rect 3451 37949 3495 38007
rect 3750 39198 3794 39242
rect 3750 39134 3794 39178
rect 4992 39135 5044 39187
rect 5034 39038 5060 39096
rect 16401 39359 16445 39417
rect 16465 39998 16509 40056
rect 5213 39038 5239 39096
rect 14721 39038 14747 39096
rect 3750 38798 3794 38842
rect 3750 38734 3794 38778
rect 4992 38735 5044 38787
rect 5034 38638 5060 38696
rect 16166 39198 16210 39242
rect 14916 39135 14968 39187
rect 16166 39134 16210 39178
rect 14900 39038 14926 39096
rect 5213 38638 5239 38696
rect 14721 38638 14747 38696
rect 16166 38798 16210 38842
rect 14916 38735 14968 38787
rect 16166 38734 16210 38778
rect 14900 38638 14926 38696
rect 5141 38560 5167 38618
rect 5320 38560 5346 38618
rect 14614 38560 14640 38618
rect 14793 38560 14819 38618
rect 3750 38398 3794 38442
rect 3750 38334 3794 38378
rect 4992 38335 5044 38387
rect 5034 38238 5060 38296
rect 5213 38238 5239 38296
rect 14721 38238 14747 38296
rect 3387 37859 3431 37917
rect 3323 36449 3367 36507
rect 3750 37998 3794 38042
rect 3750 37934 3794 37978
rect 4992 37935 5044 37987
rect 5034 37838 5060 37896
rect 16166 38398 16210 38442
rect 14916 38335 14968 38387
rect 16166 38334 16210 38378
rect 14900 38238 14926 38296
rect 5213 37838 5239 37896
rect 14721 37838 14747 37896
rect 16166 37998 16210 38042
rect 14916 37935 14968 37987
rect 16166 37934 16210 37978
rect 14900 37838 14926 37896
rect 5141 37760 5167 37818
rect 5320 37760 5346 37818
rect 14614 37760 14640 37818
rect 14793 37760 14819 37818
rect 16465 37949 16509 38007
rect 16529 39934 16573 39992
rect 16529 37859 16573 37917
rect 16593 39598 16637 39656
rect 3750 37598 3794 37642
rect 3750 37534 3794 37578
rect 4992 37535 5044 37587
rect 5034 37438 5060 37496
rect 5213 37438 5239 37496
rect 14721 37438 14747 37496
rect 3750 37198 3794 37242
rect 3750 37134 3794 37178
rect 4992 37135 5044 37187
rect 5034 37038 5060 37096
rect 16166 37598 16210 37642
rect 14916 37535 14968 37587
rect 16166 37534 16210 37578
rect 14900 37438 14926 37496
rect 5213 37038 5239 37096
rect 14721 37038 14747 37096
rect 16166 37198 16210 37242
rect 14916 37135 14968 37187
rect 16166 37134 16210 37178
rect 14900 37038 14926 37096
rect 5141 36960 5167 37018
rect 5320 36960 5346 37018
rect 14614 36960 14640 37018
rect 14793 36960 14819 37018
rect 3750 36798 3794 36842
rect 3750 36734 3794 36778
rect 4992 36735 5044 36787
rect 5034 36638 5060 36696
rect 5213 36638 5239 36696
rect 14721 36638 14747 36696
rect 3259 36359 3303 36417
rect 3195 34949 3239 35007
rect 3750 36398 3794 36442
rect 3750 36334 3794 36378
rect 4992 36335 5044 36387
rect 5034 36238 5060 36296
rect 16166 36798 16210 36842
rect 14916 36735 14968 36787
rect 16166 36734 16210 36778
rect 14900 36638 14926 36696
rect 5213 36238 5239 36296
rect 14721 36238 14747 36296
rect 16166 36398 16210 36442
rect 14916 36335 14968 36387
rect 16166 36334 16210 36378
rect 14900 36238 14926 36296
rect 5141 36160 5167 36218
rect 5320 36160 5346 36218
rect 14614 36160 14640 36218
rect 14793 36160 14819 36218
rect 16593 36449 16637 36507
rect 16657 39534 16701 39592
rect 16657 36359 16701 36417
rect 16721 39198 16765 39256
rect 3750 35998 3794 36042
rect 3750 35934 3794 35978
rect 4992 35935 5044 35987
rect 5034 35838 5060 35896
rect 5213 35838 5239 35896
rect 14721 35838 14747 35896
rect 3750 35598 3794 35642
rect 3750 35534 3794 35578
rect 4992 35535 5044 35587
rect 5034 35438 5060 35496
rect 16166 35998 16210 36042
rect 14916 35935 14968 35987
rect 16166 35934 16210 35978
rect 14900 35838 14926 35896
rect 5213 35438 5239 35496
rect 14721 35438 14747 35496
rect 16166 35598 16210 35642
rect 14916 35535 14968 35587
rect 16166 35534 16210 35578
rect 14900 35438 14926 35496
rect 5141 35360 5167 35418
rect 5320 35360 5346 35418
rect 14614 35360 14640 35418
rect 14793 35360 14819 35418
rect 3750 35198 3794 35242
rect 3750 35134 3794 35178
rect 4992 35135 5044 35187
rect 5034 35038 5060 35096
rect 5213 35038 5239 35096
rect 14721 35038 14747 35096
rect 3131 34859 3175 34917
rect 3067 33449 3111 33507
rect 3750 34798 3794 34842
rect 3750 34734 3794 34778
rect 4992 34735 5044 34787
rect 5034 34638 5060 34696
rect 16166 35198 16210 35242
rect 14916 35135 14968 35187
rect 16166 35134 16210 35178
rect 14900 35038 14926 35096
rect 16721 34949 16765 35007
rect 16785 39134 16829 39192
rect 5213 34638 5239 34696
rect 14721 34638 14747 34696
rect 16166 34798 16210 34842
rect 14916 34735 14968 34787
rect 16166 34734 16210 34778
rect 14900 34638 14926 34696
rect 5141 34560 5167 34618
rect 5320 34560 5346 34618
rect 14614 34560 14640 34618
rect 14793 34560 14819 34618
rect 16785 34859 16829 34917
rect 16849 38798 16893 38856
rect 3750 34398 3794 34442
rect 3750 34334 3794 34378
rect 4992 34335 5044 34387
rect 5034 34238 5060 34296
rect 5213 34238 5239 34296
rect 14721 34238 14747 34296
rect 3750 33998 3794 34042
rect 3750 33934 3794 33978
rect 4992 33935 5044 33987
rect 5034 33838 5060 33896
rect 16166 34398 16210 34442
rect 14916 34335 14968 34387
rect 16166 34334 16210 34378
rect 14900 34238 14926 34296
rect 5213 33838 5239 33896
rect 14721 33838 14747 33896
rect 16166 33998 16210 34042
rect 14916 33935 14968 33987
rect 16166 33934 16210 33978
rect 14900 33838 14926 33896
rect 5141 33760 5167 33818
rect 5320 33760 5346 33818
rect 14614 33760 14640 33818
rect 14793 33760 14819 33818
rect 3003 33359 3047 33417
rect 3750 33598 3794 33642
rect 3750 33534 3794 33578
rect 4992 33535 5044 33587
rect 5034 33438 5060 33496
rect 5213 33438 5239 33496
rect 14721 33438 14747 33496
rect 2939 31949 2983 32007
rect 3750 33198 3794 33242
rect 3750 33134 3794 33178
rect 4992 33135 5044 33187
rect 5034 33038 5060 33096
rect 16166 33598 16210 33642
rect 14916 33535 14968 33587
rect 16166 33534 16210 33578
rect 14900 33438 14926 33496
rect 16849 33449 16893 33507
rect 16913 38734 16957 38792
rect 16913 33359 16957 33417
rect 16977 38398 17021 38456
rect 5213 33038 5239 33096
rect 14721 33038 14747 33096
rect 16166 33198 16210 33242
rect 14916 33135 14968 33187
rect 16166 33134 16210 33178
rect 14900 33038 14926 33096
rect 5141 32960 5167 33018
rect 5320 32960 5346 33018
rect 14614 32960 14640 33018
rect 14793 32960 14819 33018
rect 3750 32798 3794 32842
rect 3750 32734 3794 32778
rect 4992 32735 5044 32787
rect 5034 32638 5060 32696
rect 5213 32638 5239 32696
rect 14721 32638 14747 32696
rect 3750 32398 3794 32442
rect 3750 32334 3794 32378
rect 4992 32335 5044 32387
rect 5034 32238 5060 32296
rect 16166 32798 16210 32842
rect 14916 32735 14968 32787
rect 16166 32734 16210 32778
rect 14900 32638 14926 32696
rect 5213 32238 5239 32296
rect 14721 32238 14747 32296
rect 16166 32398 16210 32442
rect 14916 32335 14968 32387
rect 16166 32334 16210 32378
rect 14900 32238 14926 32296
rect 5141 32160 5167 32218
rect 5320 32160 5346 32218
rect 14614 32160 14640 32218
rect 14793 32160 14819 32218
rect 2875 31859 2919 31917
rect 2811 30449 2855 30507
rect 3750 31998 3794 32042
rect 3750 31934 3794 31978
rect 4992 31935 5044 31987
rect 5034 31838 5060 31896
rect 5213 31838 5239 31896
rect 14721 31838 14747 31896
rect 3750 31598 3794 31642
rect 3750 31534 3794 31578
rect 4992 31535 5044 31587
rect 5034 31438 5060 31496
rect 16166 31998 16210 32042
rect 14916 31935 14968 31987
rect 16166 31934 16210 31978
rect 14900 31838 14926 31896
rect 16977 31949 17021 32007
rect 17041 38334 17085 38392
rect 17041 31859 17085 31917
rect 17105 38097 17149 38155
rect 5213 31438 5239 31496
rect 14721 31438 14747 31496
rect 16166 31598 16210 31642
rect 14916 31535 14968 31587
rect 16166 31534 16210 31578
rect 14900 31438 14926 31496
rect 5141 31360 5167 31418
rect 5320 31360 5346 31418
rect 14614 31360 14640 31418
rect 14793 31360 14819 31418
rect 3750 31198 3794 31242
rect 3750 31134 3794 31178
rect 4992 31135 5044 31187
rect 5034 31038 5060 31096
rect 5213 31038 5239 31096
rect 14721 31038 14747 31096
rect 3750 30798 3794 30842
rect 3750 30734 3794 30778
rect 4992 30735 5044 30787
rect 5034 30638 5060 30696
rect 16166 31198 16210 31242
rect 14916 31135 14968 31187
rect 16166 31134 16210 31178
rect 14900 31038 14926 31096
rect 5213 30638 5239 30696
rect 14721 30638 14747 30696
rect 16166 30798 16210 30842
rect 14916 30735 14968 30787
rect 16166 30734 16210 30778
rect 14900 30638 14926 30696
rect 5141 30560 5167 30618
rect 5320 30560 5346 30618
rect 14614 30560 14640 30618
rect 14793 30560 14819 30618
rect 2747 30359 2791 30417
rect 2683 28949 2727 29007
rect 3750 30398 3794 30442
rect 3750 30334 3794 30378
rect 4992 30335 5044 30387
rect 5034 30238 5060 30296
rect 5213 30238 5239 30296
rect 14721 30238 14747 30296
rect 3750 29998 3794 30042
rect 3750 29934 3794 29978
rect 4992 29935 5044 29987
rect 5034 29838 5060 29896
rect 16166 30398 16210 30442
rect 14916 30335 14968 30387
rect 16166 30334 16210 30378
rect 14900 30238 14926 30296
rect 17105 30449 17149 30507
rect 17169 38033 17213 38091
rect 17169 30359 17213 30417
rect 17233 37598 17277 37656
rect 5213 29838 5239 29896
rect 14721 29838 14747 29896
rect 16166 29998 16210 30042
rect 14916 29935 14968 29987
rect 16166 29934 16210 29978
rect 14900 29838 14926 29896
rect 5141 29760 5167 29818
rect 5320 29760 5346 29818
rect 14614 29760 14640 29818
rect 14793 29760 14819 29818
rect 3750 29598 3794 29642
rect 3750 29534 3794 29578
rect 4992 29535 5044 29587
rect 5034 29438 5060 29496
rect 5213 29438 5239 29496
rect 14721 29438 14747 29496
rect 16166 29598 16210 29642
rect 14916 29535 14968 29587
rect 16166 29534 16210 29578
rect 14900 29438 14926 29496
rect 3750 29198 3794 29242
rect 3750 29134 3794 29178
rect 4992 29135 5044 29187
rect 5034 29038 5060 29096
rect 5213 29038 5239 29096
rect 14721 29038 14747 29096
rect 16166 29198 16210 29242
rect 14916 29135 14968 29187
rect 16166 29134 16210 29178
rect 14900 29038 14926 29096
rect 2619 28859 2663 28917
rect 5175 28908 5815 28997
rect 14145 28908 14785 28997
rect 17233 28949 17277 29007
rect 17297 37534 17341 37592
rect 17297 28859 17341 28917
rect 17361 37198 17405 37256
rect 2555 27449 2599 27507
rect 17361 27449 17405 27507
rect 17425 37134 17469 37192
rect 2491 27359 2535 27417
rect 17425 27359 17469 27417
rect 17489 36798 17533 36856
rect 2427 25949 2471 26007
rect 17489 25949 17533 26007
rect 17553 36734 17597 36792
rect 2363 25859 2407 25917
rect 17553 25859 17597 25917
rect 17617 36597 17661 36655
rect 2299 24449 2343 24507
rect 17617 24449 17661 24507
rect 17681 36533 17725 36591
rect 2235 24359 2279 24417
rect 17681 24359 17725 24417
rect 17745 35998 17789 36056
rect 2171 22949 2215 23007
rect 17745 22949 17789 23007
rect 17809 35934 17853 35992
rect 2107 22859 2151 22917
rect 17809 22859 17853 22917
rect 17873 35598 17917 35656
rect 2043 21449 2087 21507
rect 17873 21449 17917 21507
rect 17937 35534 17981 35592
rect 1979 21359 2023 21417
rect 17937 21359 17981 21417
rect 18001 35198 18045 35256
rect 1915 19949 1959 20007
rect 18001 19949 18045 20007
rect 18065 35134 18109 35192
rect 1851 19859 1895 19917
rect 18065 19859 18109 19917
rect 18129 34795 18173 34853
rect 1787 18449 1831 18507
rect 18129 18449 18173 18507
rect 18193 34731 18237 34789
rect 1723 18359 1767 18417
rect 18193 18359 18237 18417
rect 18257 34398 18301 34456
rect 1659 16949 1703 17007
rect 18257 16949 18301 17007
rect 18321 34334 18365 34392
rect 1595 16859 1639 16917
rect 18321 16859 18365 16917
rect 18385 33998 18429 34056
rect 1531 15449 1575 15507
rect 18385 15449 18429 15507
rect 18449 33934 18493 33992
rect 1467 15359 1511 15417
rect 18449 15359 18493 15417
rect 18513 33598 18557 33656
rect 1403 13949 1447 14007
rect 18513 13949 18557 14007
rect 18577 33534 18621 33592
rect 1339 13859 1383 13917
rect 18577 13859 18621 13917
rect 18641 33198 18685 33256
rect 1275 12449 1319 12507
rect 18641 12449 18685 12507
rect 18705 33134 18749 33192
rect 1211 12359 1255 12417
rect 18705 12359 18749 12417
rect 18769 32798 18813 32856
rect 1147 10949 1191 11007
rect 18769 10949 18813 11007
rect 18833 32734 18877 32792
rect 1083 10859 1127 10917
rect 18833 10859 18877 10917
rect 18897 32398 18941 32456
rect 1019 9449 1063 9507
rect 18897 9449 18941 9507
rect 18961 32334 19005 32392
rect 955 9359 999 9417
rect 18961 9359 19005 9417
rect 19025 32091 19069 32149
rect 891 7949 935 8007
rect 19025 7949 19069 8007
rect 19089 32027 19133 32085
rect 827 7859 871 7917
rect 19089 7859 19133 7917
rect 19153 31598 19197 31656
rect 763 6449 807 6507
rect 19153 6449 19197 6507
rect 19217 31534 19261 31592
rect 699 6359 743 6417
rect 19217 6359 19261 6417
rect 19281 31198 19325 31256
rect 12871 6107 12965 6201
rect 12871 5483 12965 5577
rect 13009 5939 13103 6033
rect 13009 5483 13103 5577
rect 13147 5771 13241 5865
rect 13147 5483 13241 5577
rect 13285 5603 13379 5697
rect 13285 5483 13379 5577
rect 635 4949 679 5007
rect 19281 4949 19325 5007
rect 19345 31134 19389 31192
rect 571 4859 615 4917
rect 19345 4859 19389 4917
rect 19409 30798 19453 30856
rect 507 3449 551 3507
rect 19409 3449 19453 3507
rect 19473 30734 19517 30792
rect 443 3359 487 3417
rect 19473 3359 19517 3417
rect 19537 30597 19581 30655
rect 379 1949 423 2007
rect 6814 2130 6866 2156
rect 7614 2130 7666 2156
rect 8414 2130 8466 2156
rect 9214 2130 9266 2156
rect 10014 2130 10066 2156
rect 10814 2130 10866 2156
rect 11614 2130 11666 2156
rect 6086 2023 6138 2049
rect 6486 2023 6538 2049
rect 6886 2023 6938 2049
rect 7286 2023 7338 2049
rect 7686 2023 7738 2049
rect 8086 2023 8138 2049
rect 8486 2023 8538 2049
rect 8886 2023 8938 2049
rect 9286 2023 9338 2049
rect 9686 2023 9738 2049
rect 10086 2023 10138 2049
rect 10486 2023 10538 2049
rect 10886 2023 10938 2049
rect 11286 2023 11338 2049
rect 11686 2023 11738 2049
rect 12086 2023 12138 2049
rect 6814 1951 6866 1977
rect 7614 1951 7666 1977
rect 8414 1951 8466 1977
rect 9214 1951 9266 1977
rect 10014 1951 10066 1977
rect 10814 1951 10866 1977
rect 11614 1951 11666 1977
rect 315 1859 359 1917
rect 12443 1903 12517 1977
rect 19537 1949 19581 2007
rect 19601 30533 19645 30591
rect 6086 1844 6138 1870
rect 6486 1844 6538 1870
rect 6886 1844 6938 1870
rect 7286 1844 7338 1870
rect 7686 1844 7738 1870
rect 8086 1844 8138 1870
rect 8486 1844 8538 1870
rect 8886 1844 8938 1870
rect 9286 1844 9338 1870
rect 9686 1844 9738 1870
rect 10086 1844 10138 1870
rect 10486 1844 10538 1870
rect 10886 1844 10938 1870
rect 11286 1844 11338 1870
rect 11686 1844 11738 1870
rect 12086 1844 12138 1870
rect 19601 1859 19645 1917
rect 19665 29998 19709 30056
rect 251 449 295 507
rect 187 359 231 417
rect -18215 -75 -18145 -5
rect -16215 -75 -16145 -5
rect -14215 -75 -14145 -5
rect -12215 -75 -12145 -5
rect -10215 -75 -10145 -5
rect -8215 -75 -8145 -5
rect -6215 -75 -6145 -5
rect -4215 -75 -4145 -5
rect -2215 -75 -2145 -5
rect -215 -75 -145 -5
rect -18265 -1010 -18239 -984
rect -16265 -918 -16239 -892
rect -18011 -964 -17985 -938
rect -14265 -826 -14239 -800
rect -16011 -872 -15985 -846
rect -12265 -734 -12239 -708
rect -14011 -780 -13985 -754
rect -10265 -642 -10239 -616
rect -12011 -688 -11985 -662
rect -8265 -550 -8239 -524
rect -10011 -596 -9985 -570
rect -6265 -458 -6239 -432
rect -8011 -504 -7985 -478
rect -4265 -366 -4239 -340
rect -6011 -412 -5985 -386
rect -2265 -274 -2239 -248
rect -4011 -320 -3985 -294
rect -265 -182 -239 -156
rect -2011 -228 -1985 -202
rect -11 -136 15 -110
rect 19665 449 19709 507
rect 19729 29934 19773 29992
rect 19729 359 19773 417
rect 20105 -75 20175 -5
rect 22105 -75 22175 -5
rect 24105 -75 24175 -5
rect 26105 -75 26175 -5
rect 28105 -75 28175 -5
rect 30105 -75 30175 -5
rect 32105 -75 32175 -5
rect 34105 -75 34175 -5
rect 36105 -75 36175 -5
rect 38105 -75 38175 -5
rect 12250 -136 12276 -110
rect 19944 -136 19970 -110
rect 12196 -182 12222 -156
rect 11850 -228 11876 -202
rect 11796 -274 11822 -248
rect 11450 -320 11476 -294
rect 11396 -366 11422 -340
rect 11050 -412 11076 -386
rect 10996 -458 11022 -432
rect 10650 -504 10676 -478
rect 10596 -550 10622 -524
rect 10250 -596 10276 -570
rect 10196 -642 10222 -616
rect 9850 -688 9876 -662
rect 9796 -734 9822 -708
rect 9450 -780 9476 -754
rect 9396 -826 9422 -800
rect 9050 -872 9076 -846
rect 8996 -918 9022 -892
rect 8650 -964 8676 -938
rect 8596 -1010 8622 -984
rect 20198 -182 20224 -156
rect 21944 -228 21970 -202
rect 22198 -274 22224 -248
rect 23944 -320 23970 -294
rect 24198 -366 24224 -340
rect 25944 -412 25970 -386
rect 26198 -458 26224 -432
rect 27944 -504 27970 -478
rect 28198 -550 28224 -524
rect 29944 -596 29970 -570
rect 30198 -642 30224 -616
rect 31944 -688 31970 -662
rect 32198 -734 32224 -708
rect 33944 -780 33970 -754
rect 34198 -826 34224 -800
rect 35944 -872 35970 -846
rect 36198 -918 36224 -892
rect 37944 -964 37970 -938
rect 38198 -1010 38224 -984
<< metal2 >>
rect 3256 44021 3306 44024
rect 3256 44010 3259 44021
rect 40 43963 3259 44010
rect 3303 43963 3306 44021
rect 40 43960 3306 43963
rect 16654 44021 16704 44024
rect 16654 43963 16657 44021
rect 16701 44010 16704 44021
rect 16701 43963 19920 44010
rect 16654 43960 19920 43963
rect 3320 43931 3370 43934
rect 3320 43920 3323 43931
rect 40 43873 3323 43920
rect 3367 43873 3370 43931
rect 40 43870 3370 43873
rect 16590 43931 16640 43934
rect 16590 43873 16593 43931
rect 16637 43920 16640 43931
rect 16637 43873 19920 43920
rect 16590 43870 19920 43873
rect 8770 42867 11190 42872
rect 8770 42777 10923 42867
rect 11113 42777 11190 42867
rect 8770 42772 11190 42777
rect 8770 42729 11190 42734
rect 8770 42639 10655 42729
rect 10845 42639 11190 42729
rect 8770 42634 11190 42639
rect 8770 42591 11190 42596
rect 3384 42521 3434 42524
rect 3384 42510 3387 42521
rect 40 42463 3387 42510
rect 3431 42463 3434 42521
rect 8770 42501 10387 42591
rect 10577 42501 11190 42591
rect 8770 42496 11190 42501
rect 16526 42521 16576 42524
rect 40 42460 3434 42463
rect 16526 42463 16529 42521
rect 16573 42510 16576 42521
rect 16573 42463 19920 42510
rect 16526 42460 19920 42463
rect 8770 42453 11190 42458
rect 3448 42431 3498 42434
rect 3448 42420 3451 42431
rect 40 42373 3451 42420
rect 3495 42373 3498 42431
rect 40 42370 3498 42373
rect 8770 42363 10119 42453
rect 10309 42363 11190 42453
rect 16462 42431 16512 42434
rect 16462 42373 16465 42431
rect 16509 42420 16512 42431
rect 16509 42373 19920 42420
rect 16462 42370 19920 42373
rect 8770 42358 11190 42363
rect 8770 42315 11190 42320
rect 8770 42225 9851 42315
rect 10041 42225 11190 42315
rect 8770 42220 11190 42225
rect 5087 41793 5090 41871
rect 5170 41793 5320 41871
rect 14640 41793 14790 41871
rect 14870 41793 14873 41871
rect 3256 41642 3797 41645
rect 3256 41584 3259 41642
rect 3303 41598 3750 41642
rect 3794 41598 3797 41642
rect 3303 41595 3797 41598
rect 16163 41642 16704 41645
rect 16163 41598 16166 41642
rect 16210 41598 16657 41642
rect 16163 41595 16657 41598
rect 3303 41584 3306 41595
rect 3256 41581 3306 41584
rect 4989 41587 5190 41590
rect 3320 41578 3797 41581
rect 3320 41520 3323 41578
rect 3367 41534 3750 41578
rect 3794 41534 3797 41578
rect 3367 41531 3797 41534
rect 4989 41535 4992 41587
rect 5044 41535 5190 41587
rect 4989 41532 5190 41535
rect 14770 41587 14971 41590
rect 14770 41535 14916 41587
rect 14968 41535 14971 41587
rect 16654 41584 16657 41595
rect 16701 41584 16704 41642
rect 16654 41581 16704 41584
rect 14770 41532 14971 41535
rect 16163 41578 16640 41581
rect 16163 41534 16166 41578
rect 16210 41534 16593 41578
rect 16163 41531 16593 41534
rect 3367 41520 3370 41531
rect 3320 41517 3370 41520
rect 16590 41520 16593 41531
rect 16637 41520 16640 41578
rect 16590 41517 16640 41520
rect 5031 41496 5242 41499
rect 5031 41438 5034 41496
rect 5060 41438 5213 41496
rect 5239 41438 5242 41496
rect 5031 41435 5242 41438
rect 14718 41496 14929 41499
rect 14718 41438 14721 41496
rect 14747 41438 14900 41496
rect 14926 41438 14929 41496
rect 14718 41435 14929 41438
rect 3384 41242 3797 41245
rect 3384 41184 3387 41242
rect 3431 41198 3750 41242
rect 3794 41198 3797 41242
rect 3431 41195 3797 41198
rect 16163 41242 16576 41245
rect 16163 41198 16166 41242
rect 16210 41198 16529 41242
rect 16163 41195 16529 41198
rect 3431 41184 3434 41195
rect 3384 41181 3434 41184
rect 4989 41187 5190 41190
rect 3448 41178 3797 41181
rect 3448 41120 3451 41178
rect 3495 41134 3750 41178
rect 3794 41134 3797 41178
rect 3495 41131 3797 41134
rect 4989 41135 4992 41187
rect 5044 41135 5190 41187
rect 4989 41132 5190 41135
rect 14770 41187 14971 41190
rect 14770 41135 14916 41187
rect 14968 41135 14971 41187
rect 16526 41184 16529 41195
rect 16573 41184 16576 41242
rect 16526 41181 16576 41184
rect 14770 41132 14971 41135
rect 16163 41178 16512 41181
rect 16163 41134 16166 41178
rect 16210 41134 16465 41178
rect 16163 41131 16465 41134
rect 3495 41120 3498 41131
rect 3448 41117 3498 41120
rect 16462 41120 16465 41131
rect 16509 41120 16512 41178
rect 16462 41117 16512 41120
rect 5031 41096 5242 41099
rect 5031 41038 5034 41096
rect 5060 41038 5213 41096
rect 5239 41038 5242 41096
rect 5031 41035 5242 41038
rect 14718 41096 14929 41099
rect 14718 41038 14721 41096
rect 14747 41038 14900 41096
rect 14926 41038 14929 41096
rect 14718 41035 14929 41038
rect 3512 41021 3562 41024
rect 16398 41021 16448 41024
rect 3512 41010 3515 41021
rect 40 40963 3515 41010
rect 3559 40963 3562 41021
rect 40 40960 3562 40963
rect 5138 41018 5349 41021
rect 5138 40960 5141 41018
rect 5167 40960 5320 41018
rect 5346 40960 5349 41018
rect 5138 40957 5349 40960
rect 14611 41018 14822 41021
rect 14611 40960 14614 41018
rect 14640 40960 14793 41018
rect 14819 40960 14822 41018
rect 16398 40963 16401 41021
rect 16445 41010 16448 41021
rect 16445 40963 19920 41010
rect 16398 40960 19920 40963
rect 14611 40957 14822 40960
rect 3576 40931 3626 40934
rect 3576 40920 3579 40931
rect 40 40873 3579 40920
rect 3623 40873 3626 40931
rect 40 40870 3626 40873
rect 16334 40931 16384 40934
rect 16334 40873 16337 40931
rect 16381 40920 16384 40931
rect 16381 40873 19920 40920
rect 16334 40870 19920 40873
rect 3512 40842 3797 40845
rect 3512 40784 3515 40842
rect 3559 40798 3750 40842
rect 3794 40798 3797 40842
rect 3559 40795 3797 40798
rect 16163 40842 16448 40845
rect 16163 40798 16166 40842
rect 16210 40798 16401 40842
rect 16163 40795 16401 40798
rect 3559 40784 3562 40795
rect 3512 40781 3562 40784
rect 4989 40787 5190 40790
rect 3576 40778 3797 40781
rect 3576 40720 3579 40778
rect 3623 40734 3750 40778
rect 3794 40734 3797 40778
rect 3623 40731 3797 40734
rect 4989 40735 4992 40787
rect 5044 40735 5190 40787
rect 4989 40732 5190 40735
rect 14770 40787 14971 40790
rect 14770 40735 14916 40787
rect 14968 40735 14971 40787
rect 16398 40784 16401 40795
rect 16445 40784 16448 40842
rect 16398 40781 16448 40784
rect 14770 40732 14971 40735
rect 16163 40778 16384 40781
rect 16163 40734 16166 40778
rect 16210 40734 16337 40778
rect 16163 40731 16337 40734
rect 3623 40720 3626 40731
rect 3576 40717 3626 40720
rect 16334 40720 16337 40731
rect 16381 40720 16384 40778
rect 16334 40717 16384 40720
rect 5031 40696 5242 40699
rect 5031 40638 5034 40696
rect 5060 40638 5213 40696
rect 5239 40638 5242 40696
rect 5031 40635 5242 40638
rect 14718 40696 14929 40699
rect 14718 40638 14721 40696
rect 14747 40638 14900 40696
rect 14926 40638 14929 40696
rect 14718 40635 14929 40638
rect 3576 40456 3626 40459
rect 3576 40398 3579 40456
rect 3623 40445 3626 40456
rect 16334 40456 16384 40459
rect 16334 40445 16337 40456
rect 3623 40442 3797 40445
rect 3623 40398 3750 40442
rect 3794 40398 3797 40442
rect 3576 40395 3797 40398
rect 16163 40442 16337 40445
rect 16163 40398 16166 40442
rect 16210 40398 16337 40442
rect 16381 40398 16384 40456
rect 16163 40395 16384 40398
rect 3512 40392 3562 40395
rect 3512 40334 3515 40392
rect 3559 40381 3562 40392
rect 16398 40392 16448 40395
rect 4989 40387 5190 40390
rect 3559 40378 3797 40381
rect 3559 40334 3750 40378
rect 3794 40334 3797 40378
rect 3512 40331 3797 40334
rect 4989 40335 4992 40387
rect 5044 40335 5190 40387
rect 4989 40332 5190 40335
rect 14770 40387 14971 40390
rect 14770 40335 14916 40387
rect 14968 40335 14971 40387
rect 16398 40381 16401 40392
rect 14770 40332 14971 40335
rect 16163 40378 16401 40381
rect 16163 40334 16166 40378
rect 16210 40334 16401 40378
rect 16445 40334 16448 40392
rect 16163 40331 16448 40334
rect 5031 40296 5242 40299
rect 5031 40238 5034 40296
rect 5060 40238 5213 40296
rect 5239 40238 5242 40296
rect 5031 40235 5242 40238
rect 14718 40296 14929 40299
rect 14718 40238 14721 40296
rect 14747 40238 14900 40296
rect 14926 40238 14929 40296
rect 14718 40235 14929 40238
rect 5138 40218 5349 40221
rect 5138 40160 5141 40218
rect 5167 40160 5320 40218
rect 5346 40160 5349 40218
rect 5138 40157 5349 40160
rect 14611 40218 14822 40221
rect 14611 40160 14614 40218
rect 14640 40160 14793 40218
rect 14819 40160 14822 40218
rect 14611 40157 14822 40160
rect 3448 40056 3498 40059
rect 3448 39998 3451 40056
rect 3495 40045 3498 40056
rect 16462 40056 16512 40059
rect 16462 40045 16465 40056
rect 3495 40042 3797 40045
rect 3495 39998 3750 40042
rect 3794 39998 3797 40042
rect 3448 39995 3797 39998
rect 16163 40042 16465 40045
rect 16163 39998 16166 40042
rect 16210 39998 16465 40042
rect 16509 39998 16512 40056
rect 16163 39995 16512 39998
rect 3384 39992 3434 39995
rect 3384 39934 3387 39992
rect 3431 39981 3434 39992
rect 16526 39992 16576 39995
rect 4989 39987 5190 39990
rect 3431 39978 3797 39981
rect 3431 39934 3750 39978
rect 3794 39934 3797 39978
rect 3384 39931 3797 39934
rect 4989 39935 4992 39987
rect 5044 39935 5190 39987
rect 4989 39932 5190 39935
rect 14770 39987 14971 39990
rect 14770 39935 14916 39987
rect 14968 39935 14971 39987
rect 16526 39981 16529 39992
rect 14770 39932 14971 39935
rect 16163 39978 16529 39981
rect 16163 39934 16166 39978
rect 16210 39934 16529 39978
rect 16573 39934 16576 39992
rect 16163 39931 16576 39934
rect 5031 39896 5242 39899
rect 5031 39838 5034 39896
rect 5060 39838 5213 39896
rect 5239 39838 5242 39896
rect 5031 39835 5242 39838
rect 14718 39896 14929 39899
rect 14718 39838 14721 39896
rect 14747 39838 14900 39896
rect 14926 39838 14929 39896
rect 14718 39835 14929 39838
rect 3320 39656 3370 39659
rect 3320 39598 3323 39656
rect 3367 39645 3370 39656
rect 16590 39656 16640 39659
rect 16590 39645 16593 39656
rect 3367 39642 3797 39645
rect 3367 39598 3750 39642
rect 3794 39598 3797 39642
rect 3320 39595 3797 39598
rect 16163 39642 16593 39645
rect 16163 39598 16166 39642
rect 16210 39598 16593 39642
rect 16637 39598 16640 39656
rect 16163 39595 16640 39598
rect 3256 39592 3306 39595
rect 3256 39534 3259 39592
rect 3303 39581 3306 39592
rect 16654 39592 16704 39595
rect 4989 39587 5190 39590
rect 3303 39578 3797 39581
rect 3303 39534 3750 39578
rect 3794 39534 3797 39578
rect 3256 39531 3797 39534
rect 4989 39535 4992 39587
rect 5044 39535 5190 39587
rect 4989 39532 5190 39535
rect 14770 39587 14971 39590
rect 14770 39535 14916 39587
rect 14968 39535 14971 39587
rect 16654 39581 16657 39592
rect 14770 39532 14971 39535
rect 16163 39578 16657 39581
rect 16163 39534 16166 39578
rect 16210 39534 16657 39578
rect 16701 39534 16704 39592
rect 16163 39531 16704 39534
rect 40 39507 3626 39510
rect 40 39460 3579 39507
rect 3576 39449 3579 39460
rect 3623 39449 3626 39507
rect 16334 39507 19920 39510
rect 3576 39446 3626 39449
rect 5031 39496 5242 39499
rect 5031 39438 5034 39496
rect 5060 39438 5213 39496
rect 5239 39438 5242 39496
rect 5031 39435 5242 39438
rect 14718 39496 14929 39499
rect 14718 39438 14721 39496
rect 14747 39438 14900 39496
rect 14926 39438 14929 39496
rect 16334 39449 16337 39507
rect 16381 39460 19920 39507
rect 16381 39449 16384 39460
rect 16334 39446 16384 39449
rect 14718 39435 14929 39438
rect 40 39417 3562 39420
rect 40 39370 3515 39417
rect 3512 39359 3515 39370
rect 3559 39359 3562 39417
rect 3512 39356 3562 39359
rect 5138 39418 5349 39421
rect 5138 39360 5141 39418
rect 5167 39360 5320 39418
rect 5346 39360 5349 39418
rect 5138 39357 5349 39360
rect 14611 39418 14822 39421
rect 14611 39360 14614 39418
rect 14640 39360 14793 39418
rect 14819 39360 14822 39418
rect 14611 39357 14822 39360
rect 16398 39417 19920 39420
rect 16398 39359 16401 39417
rect 16445 39370 19920 39417
rect 16445 39359 16448 39370
rect 16398 39356 16448 39359
rect 3192 39256 3242 39259
rect 3192 39198 3195 39256
rect 3239 39245 3242 39256
rect 16718 39256 16768 39259
rect 16718 39245 16721 39256
rect 3239 39242 3797 39245
rect 3239 39198 3750 39242
rect 3794 39198 3797 39242
rect 3192 39195 3797 39198
rect 16163 39242 16721 39245
rect 16163 39198 16166 39242
rect 16210 39198 16721 39242
rect 16765 39198 16768 39256
rect 16163 39195 16768 39198
rect 3128 39192 3178 39195
rect 3128 39134 3131 39192
rect 3175 39181 3178 39192
rect 16782 39192 16832 39195
rect 4989 39187 5190 39190
rect 3175 39178 3797 39181
rect 3175 39134 3750 39178
rect 3794 39134 3797 39178
rect 3128 39131 3797 39134
rect 4989 39135 4992 39187
rect 5044 39135 5190 39187
rect 4989 39132 5190 39135
rect 14770 39187 14971 39190
rect 14770 39135 14916 39187
rect 14968 39135 14971 39187
rect 16782 39181 16785 39192
rect 14770 39132 14971 39135
rect 16163 39178 16785 39181
rect 16163 39134 16166 39178
rect 16210 39134 16785 39178
rect 16829 39134 16832 39192
rect 16163 39131 16832 39134
rect 5031 39096 5242 39099
rect 5031 39038 5034 39096
rect 5060 39038 5213 39096
rect 5239 39038 5242 39096
rect 5031 39035 5242 39038
rect 14718 39096 14929 39099
rect 14718 39038 14721 39096
rect 14747 39038 14900 39096
rect 14926 39038 14929 39096
rect 14718 39035 14929 39038
rect 3064 38856 3114 38859
rect 3064 38798 3067 38856
rect 3111 38845 3114 38856
rect 16846 38856 16896 38859
rect 16846 38845 16849 38856
rect 3111 38842 3797 38845
rect 3111 38798 3750 38842
rect 3794 38798 3797 38842
rect 3064 38795 3797 38798
rect 16163 38842 16849 38845
rect 16163 38798 16166 38842
rect 16210 38798 16849 38842
rect 16893 38798 16896 38856
rect 16163 38795 16896 38798
rect 3000 38792 3050 38795
rect 3000 38734 3003 38792
rect 3047 38781 3050 38792
rect 16910 38792 16960 38795
rect 4989 38787 5190 38790
rect 3047 38778 3797 38781
rect 3047 38734 3750 38778
rect 3794 38734 3797 38778
rect 3000 38731 3797 38734
rect 4989 38735 4992 38787
rect 5044 38735 5190 38787
rect 4989 38732 5190 38735
rect 14770 38787 14971 38790
rect 14770 38735 14916 38787
rect 14968 38735 14971 38787
rect 16910 38781 16913 38792
rect 14770 38732 14971 38735
rect 16163 38778 16913 38781
rect 16163 38734 16166 38778
rect 16210 38734 16913 38778
rect 16957 38734 16960 38792
rect 16163 38731 16960 38734
rect 5031 38696 5242 38699
rect 5031 38638 5034 38696
rect 5060 38638 5213 38696
rect 5239 38638 5242 38696
rect 5031 38635 5242 38638
rect 14718 38696 14929 38699
rect 14718 38638 14721 38696
rect 14747 38638 14900 38696
rect 14926 38638 14929 38696
rect 14718 38635 14929 38638
rect 5138 38618 5349 38621
rect 5138 38560 5141 38618
rect 5167 38560 5320 38618
rect 5346 38560 5349 38618
rect 5138 38557 5349 38560
rect 14611 38618 14822 38621
rect 14611 38560 14614 38618
rect 14640 38560 14793 38618
rect 14819 38560 14822 38618
rect 14611 38557 14822 38560
rect 2936 38456 2986 38459
rect 2936 38398 2939 38456
rect 2983 38445 2986 38456
rect 16974 38456 17024 38459
rect 16974 38445 16977 38456
rect 2983 38442 3797 38445
rect 2983 38398 3750 38442
rect 3794 38398 3797 38442
rect 2936 38395 3797 38398
rect 16163 38442 16977 38445
rect 16163 38398 16166 38442
rect 16210 38398 16977 38442
rect 17021 38398 17024 38456
rect 16163 38395 17024 38398
rect 2872 38392 2922 38395
rect 2872 38334 2875 38392
rect 2919 38381 2922 38392
rect 17038 38392 17088 38395
rect 4989 38387 5190 38390
rect 2919 38378 3797 38381
rect 2919 38334 3750 38378
rect 3794 38334 3797 38378
rect 2872 38331 3797 38334
rect 4989 38335 4992 38387
rect 5044 38335 5190 38387
rect 4989 38332 5190 38335
rect 14770 38387 14971 38390
rect 14770 38335 14916 38387
rect 14968 38335 14971 38387
rect 17038 38381 17041 38392
rect 14770 38332 14971 38335
rect 16163 38378 17041 38381
rect 16163 38334 16166 38378
rect 16210 38334 17041 38378
rect 17085 38334 17088 38392
rect 16163 38331 17088 38334
rect 5031 38296 5242 38299
rect 5031 38238 5034 38296
rect 5060 38238 5213 38296
rect 5239 38238 5242 38296
rect 5031 38235 5242 38238
rect 14718 38296 14929 38299
rect 14718 38238 14721 38296
rect 14747 38238 14900 38296
rect 14926 38238 14929 38296
rect 14718 38235 14929 38238
rect 2808 38155 2858 38158
rect 2808 38097 2811 38155
rect 2855 38144 2858 38155
rect 17102 38155 17152 38158
rect 17102 38144 17105 38155
rect 2855 38097 3638 38144
rect 2808 38094 3638 38097
rect 2744 38091 2794 38094
rect 2744 38033 2747 38091
rect 2791 38080 2794 38091
rect 2791 38033 3568 38080
rect 2744 38030 3568 38033
rect 40 38007 3498 38010
rect 40 37960 3451 38007
rect 3448 37949 3451 37960
rect 3495 37949 3498 38007
rect 3448 37946 3498 37949
rect 3518 37981 3568 38030
rect 3588 38045 3638 38094
rect 16322 38097 17105 38144
rect 17149 38097 17152 38155
rect 16322 38094 17152 38097
rect 16322 38045 16372 38094
rect 17166 38091 17216 38094
rect 17166 38080 17169 38091
rect 3588 38042 3797 38045
rect 3588 37998 3750 38042
rect 3794 37998 3797 38042
rect 3588 37995 3797 37998
rect 16163 38042 16372 38045
rect 16163 37998 16166 38042
rect 16210 37998 16372 38042
rect 16163 37995 16372 37998
rect 16392 38033 17169 38080
rect 17213 38033 17216 38091
rect 16392 38030 17216 38033
rect 4989 37987 5190 37990
rect 3518 37978 3797 37981
rect 3518 37934 3750 37978
rect 3794 37934 3797 37978
rect 3518 37931 3797 37934
rect 4989 37935 4992 37987
rect 5044 37935 5190 37987
rect 4989 37932 5190 37935
rect 14770 37987 14971 37990
rect 14770 37935 14916 37987
rect 14968 37935 14971 37987
rect 16392 37981 16442 38030
rect 14770 37932 14971 37935
rect 16163 37978 16442 37981
rect 16163 37934 16166 37978
rect 16210 37934 16442 37978
rect 16462 38007 19920 38010
rect 16462 37949 16465 38007
rect 16509 37960 19920 38007
rect 16509 37949 16512 37960
rect 16462 37946 16512 37949
rect 16163 37931 16442 37934
rect 40 37917 3434 37920
rect 40 37870 3387 37917
rect 3384 37859 3387 37870
rect 3431 37859 3434 37917
rect 16526 37917 19920 37920
rect 3384 37856 3434 37859
rect 5031 37896 5242 37899
rect 5031 37838 5034 37896
rect 5060 37838 5213 37896
rect 5239 37838 5242 37896
rect 5031 37835 5242 37838
rect 14718 37896 14929 37899
rect 14718 37838 14721 37896
rect 14747 37838 14900 37896
rect 14926 37838 14929 37896
rect 16526 37859 16529 37917
rect 16573 37870 19920 37917
rect 16573 37859 16576 37870
rect 16526 37856 16576 37859
rect 14718 37835 14929 37838
rect 5138 37818 5349 37821
rect 5138 37760 5141 37818
rect 5167 37760 5320 37818
rect 5346 37760 5349 37818
rect 5138 37757 5349 37760
rect 14611 37818 14822 37821
rect 14611 37760 14614 37818
rect 14640 37760 14793 37818
rect 14819 37760 14822 37818
rect 14611 37757 14822 37760
rect 2680 37656 2730 37659
rect 2680 37598 2683 37656
rect 2727 37645 2730 37656
rect 17230 37656 17280 37659
rect 17230 37645 17233 37656
rect 2727 37642 3797 37645
rect 2727 37598 3750 37642
rect 3794 37598 3797 37642
rect 2680 37595 3797 37598
rect 16163 37642 17233 37645
rect 16163 37598 16166 37642
rect 16210 37598 17233 37642
rect 17277 37598 17280 37656
rect 16163 37595 17280 37598
rect 2616 37592 2666 37595
rect 2616 37534 2619 37592
rect 2663 37581 2666 37592
rect 17294 37592 17344 37595
rect 4989 37587 5190 37590
rect 2663 37578 3797 37581
rect 2663 37534 3750 37578
rect 3794 37534 3797 37578
rect 2616 37531 3797 37534
rect 4989 37535 4992 37587
rect 5044 37535 5190 37587
rect 4989 37532 5190 37535
rect 14770 37587 14971 37590
rect 14770 37535 14916 37587
rect 14968 37535 14971 37587
rect 17294 37581 17297 37592
rect 14770 37532 14971 37535
rect 16163 37578 17297 37581
rect 16163 37534 16166 37578
rect 16210 37534 17297 37578
rect 17341 37534 17344 37592
rect 16163 37531 17344 37534
rect 5031 37496 5242 37499
rect 5031 37438 5034 37496
rect 5060 37438 5213 37496
rect 5239 37438 5242 37496
rect 5031 37435 5242 37438
rect 14718 37496 14929 37499
rect 14718 37438 14721 37496
rect 14747 37438 14900 37496
rect 14926 37438 14929 37496
rect 14718 37435 14929 37438
rect 2552 37256 2602 37259
rect 2552 37198 2555 37256
rect 2599 37245 2602 37256
rect 17358 37256 17408 37259
rect 17358 37245 17361 37256
rect 2599 37242 3797 37245
rect 2599 37198 3750 37242
rect 3794 37198 3797 37242
rect 2552 37195 3797 37198
rect 16163 37242 17361 37245
rect 16163 37198 16166 37242
rect 16210 37198 17361 37242
rect 17405 37198 17408 37256
rect 16163 37195 17408 37198
rect 2488 37192 2538 37195
rect 2488 37134 2491 37192
rect 2535 37181 2538 37192
rect 17422 37192 17472 37195
rect 4989 37187 5190 37190
rect 2535 37178 3797 37181
rect 2535 37134 3750 37178
rect 3794 37134 3797 37178
rect 2488 37131 3797 37134
rect 4989 37135 4992 37187
rect 5044 37135 5190 37187
rect 4989 37132 5190 37135
rect 14770 37187 14971 37190
rect 14770 37135 14916 37187
rect 14968 37135 14971 37187
rect 17422 37181 17425 37192
rect 14770 37132 14971 37135
rect 16163 37178 17425 37181
rect 16163 37134 16166 37178
rect 16210 37134 17425 37178
rect 17469 37134 17472 37192
rect 16163 37131 17472 37134
rect 5031 37096 5242 37099
rect 5031 37038 5034 37096
rect 5060 37038 5213 37096
rect 5239 37038 5242 37096
rect 5031 37035 5242 37038
rect 14718 37096 14929 37099
rect 14718 37038 14721 37096
rect 14747 37038 14900 37096
rect 14926 37038 14929 37096
rect 14718 37035 14929 37038
rect 5138 37018 5349 37021
rect 5138 36960 5141 37018
rect 5167 36960 5320 37018
rect 5346 36960 5349 37018
rect 5138 36957 5349 36960
rect 14611 37018 14822 37021
rect 14611 36960 14614 37018
rect 14640 36960 14793 37018
rect 14819 36960 14822 37018
rect 14611 36957 14822 36960
rect 2424 36856 2474 36859
rect 2424 36798 2427 36856
rect 2471 36845 2474 36856
rect 17486 36856 17536 36859
rect 17486 36845 17489 36856
rect 2471 36842 3797 36845
rect 2471 36798 3750 36842
rect 3794 36798 3797 36842
rect 2424 36795 3797 36798
rect 16163 36842 17489 36845
rect 16163 36798 16166 36842
rect 16210 36798 17489 36842
rect 17533 36798 17536 36856
rect 16163 36795 17536 36798
rect 2360 36792 2410 36795
rect 2360 36734 2363 36792
rect 2407 36781 2410 36792
rect 17550 36792 17600 36795
rect 4989 36787 5190 36790
rect 2407 36778 3797 36781
rect 2407 36734 3750 36778
rect 3794 36734 3797 36778
rect 2360 36731 3797 36734
rect 4989 36735 4992 36787
rect 5044 36735 5190 36787
rect 4989 36732 5190 36735
rect 14770 36787 14971 36790
rect 14770 36735 14916 36787
rect 14968 36735 14971 36787
rect 17550 36781 17553 36792
rect 14770 36732 14971 36735
rect 16163 36778 17553 36781
rect 16163 36734 16166 36778
rect 16210 36734 17553 36778
rect 17597 36734 17600 36792
rect 16163 36731 17600 36734
rect 5031 36696 5242 36699
rect 2296 36655 2346 36658
rect 2296 36597 2299 36655
rect 2343 36644 2346 36655
rect 2343 36597 3588 36644
rect 5031 36638 5034 36696
rect 5060 36638 5213 36696
rect 5239 36638 5242 36696
rect 5031 36635 5242 36638
rect 14718 36696 14929 36699
rect 14718 36638 14721 36696
rect 14747 36638 14900 36696
rect 14926 36638 14929 36696
rect 17614 36655 17664 36658
rect 17614 36644 17617 36655
rect 14718 36635 14929 36638
rect 2296 36594 3588 36597
rect 2232 36591 2282 36594
rect 2232 36533 2235 36591
rect 2279 36580 2282 36591
rect 2279 36533 3518 36580
rect 2232 36530 3518 36533
rect 40 36507 3370 36510
rect 40 36460 3323 36507
rect 3320 36449 3323 36460
rect 3367 36449 3370 36507
rect 3320 36446 3370 36449
rect 40 36417 3306 36420
rect 40 36370 3259 36417
rect 3256 36359 3259 36370
rect 3303 36359 3306 36417
rect 3256 36356 3306 36359
rect 3468 36381 3518 36530
rect 3538 36445 3588 36594
rect 16372 36597 17617 36644
rect 17661 36597 17664 36655
rect 16372 36594 17664 36597
rect 16372 36445 16422 36594
rect 17678 36591 17728 36594
rect 17678 36580 17681 36591
rect 3538 36442 3797 36445
rect 3538 36398 3750 36442
rect 3794 36398 3797 36442
rect 3538 36395 3797 36398
rect 16163 36442 16422 36445
rect 16163 36398 16166 36442
rect 16210 36398 16422 36442
rect 16163 36395 16422 36398
rect 16442 36533 17681 36580
rect 17725 36533 17728 36591
rect 16442 36530 17728 36533
rect 4989 36387 5190 36390
rect 3468 36378 3797 36381
rect 3468 36334 3750 36378
rect 3794 36334 3797 36378
rect 3468 36331 3797 36334
rect 4989 36335 4992 36387
rect 5044 36335 5190 36387
rect 4989 36332 5190 36335
rect 14770 36387 14971 36390
rect 14770 36335 14916 36387
rect 14968 36335 14971 36387
rect 16442 36381 16492 36530
rect 16590 36507 19920 36510
rect 16590 36449 16593 36507
rect 16637 36460 19920 36507
rect 16637 36449 16640 36460
rect 16590 36446 16640 36449
rect 14770 36332 14971 36335
rect 16163 36378 16492 36381
rect 16163 36334 16166 36378
rect 16210 36334 16492 36378
rect 16654 36417 19920 36420
rect 16654 36359 16657 36417
rect 16701 36370 19920 36417
rect 16701 36359 16704 36370
rect 16654 36356 16704 36359
rect 16163 36331 16492 36334
rect 5031 36296 5242 36299
rect 5031 36238 5034 36296
rect 5060 36238 5213 36296
rect 5239 36238 5242 36296
rect 5031 36235 5242 36238
rect 14718 36296 14929 36299
rect 14718 36238 14721 36296
rect 14747 36238 14900 36296
rect 14926 36238 14929 36296
rect 14718 36235 14929 36238
rect 5138 36218 5349 36221
rect 5138 36160 5141 36218
rect 5167 36160 5320 36218
rect 5346 36160 5349 36218
rect 5138 36157 5349 36160
rect 14611 36218 14822 36221
rect 14611 36160 14614 36218
rect 14640 36160 14793 36218
rect 14819 36160 14822 36218
rect 14611 36157 14822 36160
rect 2168 36056 2218 36059
rect 2168 35998 2171 36056
rect 2215 36045 2218 36056
rect 17742 36056 17792 36059
rect 17742 36045 17745 36056
rect 2215 36042 3797 36045
rect 2215 35998 3750 36042
rect 3794 35998 3797 36042
rect 2168 35995 3797 35998
rect 16163 36042 17745 36045
rect 16163 35998 16166 36042
rect 16210 35998 17745 36042
rect 17789 35998 17792 36056
rect 16163 35995 17792 35998
rect 2104 35992 2154 35995
rect 2104 35934 2107 35992
rect 2151 35981 2154 35992
rect 17806 35992 17856 35995
rect 4989 35987 5190 35990
rect 2151 35978 3797 35981
rect 2151 35934 3750 35978
rect 3794 35934 3797 35978
rect 2104 35931 3797 35934
rect 4989 35935 4992 35987
rect 5044 35935 5190 35987
rect 4989 35932 5190 35935
rect 14770 35987 14971 35990
rect 14770 35935 14916 35987
rect 14968 35935 14971 35987
rect 17806 35981 17809 35992
rect 14770 35932 14971 35935
rect 16163 35978 17809 35981
rect 16163 35934 16166 35978
rect 16210 35934 17809 35978
rect 17853 35934 17856 35992
rect 16163 35931 17856 35934
rect 5031 35896 5242 35899
rect 5031 35838 5034 35896
rect 5060 35838 5213 35896
rect 5239 35838 5242 35896
rect 5031 35835 5242 35838
rect 14718 35896 14929 35899
rect 14718 35838 14721 35896
rect 14747 35838 14900 35896
rect 14926 35838 14929 35896
rect 14718 35835 14929 35838
rect 2040 35656 2090 35659
rect 2040 35598 2043 35656
rect 2087 35645 2090 35656
rect 17870 35656 17920 35659
rect 17870 35645 17873 35656
rect 2087 35642 3797 35645
rect 2087 35598 3750 35642
rect 3794 35598 3797 35642
rect 2040 35595 3797 35598
rect 16163 35642 17873 35645
rect 16163 35598 16166 35642
rect 16210 35598 17873 35642
rect 17917 35598 17920 35656
rect 16163 35595 17920 35598
rect 1976 35592 2026 35595
rect 1976 35534 1979 35592
rect 2023 35581 2026 35592
rect 17934 35592 17984 35595
rect 4989 35587 5190 35590
rect 2023 35578 3797 35581
rect 2023 35534 3750 35578
rect 3794 35534 3797 35578
rect 1976 35531 3797 35534
rect 4989 35535 4992 35587
rect 5044 35535 5190 35587
rect 4989 35532 5190 35535
rect 14770 35587 14971 35590
rect 14770 35535 14916 35587
rect 14968 35535 14971 35587
rect 17934 35581 17937 35592
rect 14770 35532 14971 35535
rect 16163 35578 17937 35581
rect 16163 35534 16166 35578
rect 16210 35534 17937 35578
rect 17981 35534 17984 35592
rect 16163 35531 17984 35534
rect 5031 35496 5242 35499
rect 5031 35438 5034 35496
rect 5060 35438 5213 35496
rect 5239 35438 5242 35496
rect 5031 35435 5242 35438
rect 14718 35496 14929 35499
rect 14718 35438 14721 35496
rect 14747 35438 14900 35496
rect 14926 35438 14929 35496
rect 14718 35435 14929 35438
rect 5138 35418 5349 35421
rect 5138 35360 5141 35418
rect 5167 35360 5320 35418
rect 5346 35360 5349 35418
rect 5138 35357 5349 35360
rect 14611 35418 14822 35421
rect 14611 35360 14614 35418
rect 14640 35360 14793 35418
rect 14819 35360 14822 35418
rect 14611 35357 14822 35360
rect 1912 35256 1962 35259
rect 1912 35198 1915 35256
rect 1959 35245 1962 35256
rect 17998 35256 18048 35259
rect 17998 35245 18001 35256
rect 1959 35242 3797 35245
rect 1959 35198 3750 35242
rect 3794 35198 3797 35242
rect 1912 35195 3797 35198
rect 16163 35242 18001 35245
rect 16163 35198 16166 35242
rect 16210 35198 18001 35242
rect 18045 35198 18048 35256
rect 16163 35195 18048 35198
rect 1848 35192 1898 35195
rect 1848 35134 1851 35192
rect 1895 35181 1898 35192
rect 18062 35192 18112 35195
rect 4989 35187 5190 35190
rect 1895 35178 3797 35181
rect 1895 35134 3750 35178
rect 3794 35134 3797 35178
rect 1848 35131 3797 35134
rect 4989 35135 4992 35187
rect 5044 35135 5190 35187
rect 4989 35132 5190 35135
rect 14770 35187 14971 35190
rect 14770 35135 14916 35187
rect 14968 35135 14971 35187
rect 18062 35181 18065 35192
rect 14770 35132 14971 35135
rect 16163 35178 18065 35181
rect 16163 35134 16166 35178
rect 16210 35134 18065 35178
rect 18109 35134 18112 35192
rect 16163 35131 18112 35134
rect 5031 35096 5242 35099
rect 5031 35038 5034 35096
rect 5060 35038 5213 35096
rect 5239 35038 5242 35096
rect 5031 35035 5242 35038
rect 14718 35096 14929 35099
rect 14718 35038 14721 35096
rect 14747 35038 14900 35096
rect 14926 35038 14929 35096
rect 14718 35035 14929 35038
rect 40 35007 3242 35010
rect 40 34960 3195 35007
rect 3192 34949 3195 34960
rect 3239 34949 3242 35007
rect 3192 34946 3242 34949
rect 16718 35007 19920 35010
rect 16718 34949 16721 35007
rect 16765 34960 19920 35007
rect 16765 34949 16768 34960
rect 16718 34946 16768 34949
rect 40 34917 3178 34920
rect 40 34870 3131 34917
rect 3128 34859 3131 34870
rect 3175 34859 3178 34917
rect 3128 34856 3178 34859
rect 16782 34917 19920 34920
rect 16782 34859 16785 34917
rect 16829 34870 19920 34917
rect 16829 34859 16832 34870
rect 16782 34856 16832 34859
rect 1784 34853 1834 34856
rect 1784 34795 1787 34853
rect 1831 34842 1834 34853
rect 18126 34853 18176 34856
rect 3193 34842 3797 34845
rect 1831 34798 3750 34842
rect 3794 34798 3797 34842
rect 1831 34795 3797 34798
rect 16163 34842 16767 34845
rect 18126 34842 18129 34853
rect 16163 34798 16166 34842
rect 16210 34798 18129 34842
rect 16163 34795 18129 34798
rect 18173 34795 18176 34853
rect 1784 34792 3207 34795
rect 16753 34792 18176 34795
rect 1720 34789 1770 34792
rect 1720 34731 1723 34789
rect 1767 34778 1770 34789
rect 4989 34787 5190 34790
rect 3216 34778 3797 34781
rect 1767 34734 3750 34778
rect 3794 34734 3797 34778
rect 1767 34731 3797 34734
rect 4989 34735 4992 34787
rect 5044 34735 5190 34787
rect 4989 34732 5190 34735
rect 14770 34787 14971 34790
rect 14770 34735 14916 34787
rect 14968 34735 14971 34787
rect 18190 34789 18240 34792
rect 14770 34732 14971 34735
rect 16163 34778 16744 34781
rect 18190 34778 18193 34789
rect 16163 34734 16166 34778
rect 16210 34734 18193 34778
rect 16163 34731 18193 34734
rect 18237 34731 18240 34789
rect 1720 34728 3230 34731
rect 16730 34728 18240 34731
rect 5031 34696 5242 34699
rect 5031 34638 5034 34696
rect 5060 34638 5213 34696
rect 5239 34638 5242 34696
rect 5031 34635 5242 34638
rect 14718 34696 14929 34699
rect 14718 34638 14721 34696
rect 14747 34638 14900 34696
rect 14926 34638 14929 34696
rect 14718 34635 14929 34638
rect 5138 34618 5349 34621
rect 5138 34560 5141 34618
rect 5167 34560 5320 34618
rect 5346 34560 5349 34618
rect 5138 34557 5349 34560
rect 14611 34618 14822 34621
rect 14611 34560 14614 34618
rect 14640 34560 14793 34618
rect 14819 34560 14822 34618
rect 14611 34557 14822 34560
rect 1656 34456 1706 34459
rect 1656 34398 1659 34456
rect 1703 34445 1706 34456
rect 18254 34456 18304 34459
rect 18254 34445 18257 34456
rect 1703 34442 3797 34445
rect 1703 34398 3750 34442
rect 3794 34398 3797 34442
rect 1656 34395 3797 34398
rect 16163 34442 18257 34445
rect 16163 34398 16166 34442
rect 16210 34398 18257 34442
rect 18301 34398 18304 34456
rect 16163 34395 18304 34398
rect 1592 34392 1642 34395
rect 1592 34334 1595 34392
rect 1639 34381 1642 34392
rect 18318 34392 18368 34395
rect 4989 34387 5190 34390
rect 1639 34378 3797 34381
rect 1639 34334 3750 34378
rect 3794 34334 3797 34378
rect 1592 34331 3797 34334
rect 4989 34335 4992 34387
rect 5044 34335 5190 34387
rect 4989 34332 5190 34335
rect 14770 34387 14971 34390
rect 14770 34335 14916 34387
rect 14968 34335 14971 34387
rect 18318 34381 18321 34392
rect 14770 34332 14971 34335
rect 16163 34378 18321 34381
rect 16163 34334 16166 34378
rect 16210 34334 18321 34378
rect 18365 34334 18368 34392
rect 16163 34331 18368 34334
rect 5031 34296 5242 34299
rect 5031 34238 5034 34296
rect 5060 34238 5213 34296
rect 5239 34238 5242 34296
rect 5031 34235 5242 34238
rect 14718 34296 14929 34299
rect 14718 34238 14721 34296
rect 14747 34238 14900 34296
rect 14926 34238 14929 34296
rect 14718 34235 14929 34238
rect 1528 34056 1578 34059
rect 1528 33998 1531 34056
rect 1575 34045 1578 34056
rect 18382 34056 18432 34059
rect 18382 34045 18385 34056
rect 1575 34042 3797 34045
rect 1575 33998 3750 34042
rect 3794 33998 3797 34042
rect 1528 33995 3797 33998
rect 16163 34042 18385 34045
rect 16163 33998 16166 34042
rect 16210 33998 18385 34042
rect 18429 33998 18432 34056
rect 16163 33995 18432 33998
rect 1464 33992 1514 33995
rect 1464 33934 1467 33992
rect 1511 33981 1514 33992
rect 18446 33992 18496 33995
rect 4989 33987 5190 33990
rect 1511 33978 3797 33981
rect 1511 33934 3750 33978
rect 3794 33934 3797 33978
rect 1464 33931 3797 33934
rect 4989 33935 4992 33987
rect 5044 33935 5190 33987
rect 4989 33932 5190 33935
rect 14770 33987 14971 33990
rect 14770 33935 14916 33987
rect 14968 33935 14971 33987
rect 18446 33981 18449 33992
rect 14770 33932 14971 33935
rect 16163 33978 18449 33981
rect 16163 33934 16166 33978
rect 16210 33934 18449 33978
rect 18493 33934 18496 33992
rect 16163 33931 18496 33934
rect 5031 33896 5242 33899
rect 5031 33838 5034 33896
rect 5060 33838 5213 33896
rect 5239 33838 5242 33896
rect 5031 33835 5242 33838
rect 14718 33896 14929 33899
rect 14718 33838 14721 33896
rect 14747 33838 14900 33896
rect 14926 33838 14929 33896
rect 14718 33835 14929 33838
rect 5138 33818 5349 33821
rect 5138 33760 5141 33818
rect 5167 33760 5320 33818
rect 5346 33760 5349 33818
rect 5138 33757 5349 33760
rect 14611 33818 14822 33821
rect 14611 33760 14614 33818
rect 14640 33760 14793 33818
rect 14819 33760 14822 33818
rect 14611 33757 14822 33760
rect 1400 33656 1450 33659
rect 1400 33598 1403 33656
rect 1447 33645 1450 33656
rect 18510 33656 18560 33659
rect 18510 33645 18513 33656
rect 1447 33642 3797 33645
rect 1447 33598 3750 33642
rect 3794 33598 3797 33642
rect 1400 33595 3797 33598
rect 16163 33642 18513 33645
rect 16163 33598 16166 33642
rect 16210 33598 18513 33642
rect 18557 33598 18560 33656
rect 16163 33595 18560 33598
rect 1336 33592 1386 33595
rect 1336 33534 1339 33592
rect 1383 33581 1386 33592
rect 18574 33592 18624 33595
rect 4989 33587 5190 33590
rect 1383 33578 3797 33581
rect 1383 33534 3750 33578
rect 3794 33534 3797 33578
rect 1336 33531 3797 33534
rect 4989 33535 4992 33587
rect 5044 33535 5190 33587
rect 4989 33532 5190 33535
rect 14770 33587 14971 33590
rect 14770 33535 14916 33587
rect 14968 33535 14971 33587
rect 18574 33581 18577 33592
rect 14770 33532 14971 33535
rect 16163 33578 18577 33581
rect 16163 33534 16166 33578
rect 16210 33534 18577 33578
rect 18621 33534 18624 33592
rect 16163 33531 18624 33534
rect 40 33507 3114 33510
rect 40 33460 3067 33507
rect 3064 33449 3067 33460
rect 3111 33449 3114 33507
rect 16846 33507 19920 33510
rect 3064 33446 3114 33449
rect 5031 33496 5242 33499
rect 5031 33438 5034 33496
rect 5060 33438 5213 33496
rect 5239 33438 5242 33496
rect 5031 33435 5242 33438
rect 14718 33496 14929 33499
rect 14718 33438 14721 33496
rect 14747 33438 14900 33496
rect 14926 33438 14929 33496
rect 16846 33449 16849 33507
rect 16893 33460 19920 33507
rect 16893 33449 16896 33460
rect 16846 33446 16896 33449
rect 14718 33435 14929 33438
rect 40 33417 3050 33420
rect 40 33370 3003 33417
rect 3000 33359 3003 33370
rect 3047 33359 3050 33417
rect 3000 33356 3050 33359
rect 16910 33417 19920 33420
rect 16910 33359 16913 33417
rect 16957 33370 19920 33417
rect 16957 33359 16960 33370
rect 16910 33356 16960 33359
rect 1272 33256 1322 33259
rect 1272 33198 1275 33256
rect 1319 33245 1322 33256
rect 18638 33256 18688 33259
rect 18638 33245 18641 33256
rect 1319 33242 3797 33245
rect 1319 33198 3750 33242
rect 3794 33198 3797 33242
rect 1272 33195 3797 33198
rect 16163 33242 18641 33245
rect 16163 33198 16166 33242
rect 16210 33198 18641 33242
rect 18685 33198 18688 33256
rect 16163 33195 18688 33198
rect 1208 33192 1258 33195
rect 1208 33134 1211 33192
rect 1255 33181 1258 33192
rect 18702 33192 18752 33195
rect 4989 33187 5190 33190
rect 1255 33178 3797 33181
rect 1255 33134 3750 33178
rect 3794 33134 3797 33178
rect 1208 33131 3797 33134
rect 4989 33135 4992 33187
rect 5044 33135 5190 33187
rect 4989 33132 5190 33135
rect 14770 33187 14971 33190
rect 14770 33135 14916 33187
rect 14968 33135 14971 33187
rect 18702 33181 18705 33192
rect 14770 33132 14971 33135
rect 16163 33178 18705 33181
rect 16163 33134 16166 33178
rect 16210 33134 18705 33178
rect 18749 33134 18752 33192
rect 16163 33131 18752 33134
rect 5031 33096 5242 33099
rect 5031 33038 5034 33096
rect 5060 33038 5213 33096
rect 5239 33038 5242 33096
rect 5031 33035 5242 33038
rect 14718 33096 14929 33099
rect 14718 33038 14721 33096
rect 14747 33038 14900 33096
rect 14926 33038 14929 33096
rect 14718 33035 14929 33038
rect 5138 33018 5349 33021
rect 5138 32960 5141 33018
rect 5167 32960 5320 33018
rect 5346 32960 5349 33018
rect 5138 32957 5349 32960
rect 14611 33018 14822 33021
rect 14611 32960 14614 33018
rect 14640 32960 14793 33018
rect 14819 32960 14822 33018
rect 14611 32957 14822 32960
rect 1144 32856 1194 32859
rect 1144 32798 1147 32856
rect 1191 32845 1194 32856
rect 18766 32856 18816 32859
rect 18766 32845 18769 32856
rect 1191 32842 3797 32845
rect 1191 32798 3750 32842
rect 3794 32798 3797 32842
rect 1144 32795 3797 32798
rect 16163 32842 18769 32845
rect 16163 32798 16166 32842
rect 16210 32798 18769 32842
rect 18813 32798 18816 32856
rect 16163 32795 18816 32798
rect 1080 32792 1130 32795
rect 1080 32734 1083 32792
rect 1127 32781 1130 32792
rect 18830 32792 18880 32795
rect 4989 32787 5190 32790
rect 1127 32778 3797 32781
rect 1127 32734 3750 32778
rect 3794 32734 3797 32778
rect 1080 32731 3797 32734
rect 4989 32735 4992 32787
rect 5044 32735 5190 32787
rect 4989 32732 5190 32735
rect 14770 32787 14971 32790
rect 14770 32735 14916 32787
rect 14968 32735 14971 32787
rect 18830 32781 18833 32792
rect 14770 32732 14971 32735
rect 16163 32778 18833 32781
rect 16163 32734 16166 32778
rect 16210 32734 18833 32778
rect 18877 32734 18880 32792
rect 16163 32731 18880 32734
rect 5031 32696 5242 32699
rect 5031 32638 5034 32696
rect 5060 32638 5213 32696
rect 5239 32638 5242 32696
rect 5031 32635 5242 32638
rect 14718 32696 14929 32699
rect 14718 32638 14721 32696
rect 14747 32638 14900 32696
rect 14926 32638 14929 32696
rect 14718 32635 14929 32638
rect 1016 32456 1066 32459
rect 1016 32398 1019 32456
rect 1063 32445 1066 32456
rect 18894 32456 18944 32459
rect 18894 32445 18897 32456
rect 1063 32442 3797 32445
rect 1063 32398 3750 32442
rect 3794 32398 3797 32442
rect 1016 32395 3797 32398
rect 16163 32442 18897 32445
rect 16163 32398 16166 32442
rect 16210 32398 18897 32442
rect 18941 32398 18944 32456
rect 16163 32395 18944 32398
rect 952 32392 1002 32395
rect 952 32334 955 32392
rect 999 32381 1002 32392
rect 18958 32392 19008 32395
rect 4989 32387 5190 32390
rect 999 32378 3797 32381
rect 999 32334 3750 32378
rect 3794 32334 3797 32378
rect 952 32331 3797 32334
rect 4989 32335 4992 32387
rect 5044 32335 5190 32387
rect 4989 32332 5190 32335
rect 14770 32387 14971 32390
rect 14770 32335 14916 32387
rect 14968 32335 14971 32387
rect 18958 32381 18961 32392
rect 14770 32332 14971 32335
rect 16163 32378 18961 32381
rect 16163 32334 16166 32378
rect 16210 32334 18961 32378
rect 19005 32334 19008 32392
rect 16163 32331 19008 32334
rect 5031 32296 5242 32299
rect 5031 32238 5034 32296
rect 5060 32238 5213 32296
rect 5239 32238 5242 32296
rect 5031 32235 5242 32238
rect 14718 32296 14929 32299
rect 14718 32238 14721 32296
rect 14747 32238 14900 32296
rect 14926 32238 14929 32296
rect 14718 32235 14929 32238
rect 5138 32218 5349 32221
rect 5138 32160 5141 32218
rect 5167 32160 5320 32218
rect 5346 32160 5349 32218
rect 5138 32157 5349 32160
rect 14611 32218 14822 32221
rect 14611 32160 14614 32218
rect 14640 32160 14793 32218
rect 14819 32160 14822 32218
rect 14611 32157 14822 32160
rect 888 32149 938 32152
rect 888 32091 891 32149
rect 935 32138 938 32149
rect 19022 32149 19072 32152
rect 19022 32138 19025 32149
rect 935 32091 3588 32138
rect 888 32088 3588 32091
rect 824 32085 874 32088
rect 824 32027 827 32085
rect 871 32074 874 32085
rect 871 32027 3518 32074
rect 824 32024 3518 32027
rect 40 32007 2986 32010
rect 40 31960 2939 32007
rect 2936 31949 2939 31960
rect 2983 31949 2986 32007
rect 2936 31946 2986 31949
rect 3468 31981 3518 32024
rect 3538 32045 3588 32088
rect 16372 32091 19025 32138
rect 19069 32091 19072 32149
rect 16372 32088 19072 32091
rect 16372 32045 16422 32088
rect 19086 32085 19136 32088
rect 19086 32074 19089 32085
rect 3538 32042 3797 32045
rect 3538 31998 3750 32042
rect 3794 31998 3797 32042
rect 3538 31995 3797 31998
rect 16163 32042 16422 32045
rect 16163 31998 16166 32042
rect 16210 31998 16422 32042
rect 16163 31995 16422 31998
rect 16442 32027 19089 32074
rect 19133 32027 19136 32085
rect 16442 32024 19136 32027
rect 4989 31987 5190 31990
rect 3468 31978 3797 31981
rect 3468 31934 3750 31978
rect 3794 31934 3797 31978
rect 3468 31931 3797 31934
rect 4989 31935 4992 31987
rect 5044 31935 5190 31987
rect 4989 31932 5190 31935
rect 14770 31987 14971 31990
rect 14770 31935 14916 31987
rect 14968 31935 14971 31987
rect 16442 31981 16492 32024
rect 14770 31932 14971 31935
rect 16163 31978 16492 31981
rect 16163 31934 16166 31978
rect 16210 31934 16492 31978
rect 16974 32007 19920 32010
rect 16974 31949 16977 32007
rect 17021 31960 19920 32007
rect 17021 31949 17024 31960
rect 16974 31946 17024 31949
rect 16163 31931 16492 31934
rect 40 31917 2922 31920
rect 40 31870 2875 31917
rect 2872 31859 2875 31870
rect 2919 31859 2922 31917
rect 17038 31917 19920 31920
rect 2872 31856 2922 31859
rect 5031 31896 5242 31899
rect 5031 31838 5034 31896
rect 5060 31838 5213 31896
rect 5239 31838 5242 31896
rect 5031 31835 5242 31838
rect 14718 31896 14929 31899
rect 14718 31838 14721 31896
rect 14747 31838 14900 31896
rect 14926 31838 14929 31896
rect 17038 31859 17041 31917
rect 17085 31870 19920 31917
rect 17085 31859 17088 31870
rect 17038 31856 17088 31859
rect 14718 31835 14929 31838
rect 760 31656 810 31659
rect 760 31598 763 31656
rect 807 31645 810 31656
rect 19150 31656 19200 31659
rect 19150 31645 19153 31656
rect 807 31642 3797 31645
rect 807 31598 3750 31642
rect 3794 31598 3797 31642
rect 760 31595 3797 31598
rect 16163 31642 19153 31645
rect 16163 31598 16166 31642
rect 16210 31598 19153 31642
rect 19197 31598 19200 31656
rect 16163 31595 19200 31598
rect 696 31592 746 31595
rect 696 31534 699 31592
rect 743 31581 746 31592
rect 19214 31592 19264 31595
rect 4989 31587 5190 31590
rect 743 31578 3797 31581
rect 743 31534 3750 31578
rect 3794 31534 3797 31578
rect 696 31531 3797 31534
rect 4989 31535 4992 31587
rect 5044 31535 5190 31587
rect 4989 31532 5190 31535
rect 14770 31587 14971 31590
rect 14770 31535 14916 31587
rect 14968 31535 14971 31587
rect 19214 31581 19217 31592
rect 14770 31532 14971 31535
rect 16163 31578 19217 31581
rect 16163 31534 16166 31578
rect 16210 31534 19217 31578
rect 19261 31534 19264 31592
rect 16163 31531 19264 31534
rect 5031 31496 5242 31499
rect 5031 31438 5034 31496
rect 5060 31438 5213 31496
rect 5239 31438 5242 31496
rect 5031 31435 5242 31438
rect 14718 31496 14929 31499
rect 14718 31438 14721 31496
rect 14747 31438 14900 31496
rect 14926 31438 14929 31496
rect 14718 31435 14929 31438
rect 5138 31418 5349 31421
rect 5138 31360 5141 31418
rect 5167 31360 5320 31418
rect 5346 31360 5349 31418
rect 5138 31357 5349 31360
rect 14611 31418 14822 31421
rect 14611 31360 14614 31418
rect 14640 31360 14793 31418
rect 14819 31360 14822 31418
rect 14611 31357 14822 31360
rect 632 31256 682 31259
rect 632 31198 635 31256
rect 679 31245 682 31256
rect 19278 31256 19328 31259
rect 19278 31245 19281 31256
rect 679 31242 3797 31245
rect 679 31198 3750 31242
rect 3794 31198 3797 31242
rect 632 31195 3797 31198
rect 16163 31242 19281 31245
rect 16163 31198 16166 31242
rect 16210 31198 19281 31242
rect 19325 31198 19328 31256
rect 16163 31195 19328 31198
rect 568 31192 618 31195
rect 568 31134 571 31192
rect 615 31181 618 31192
rect 19342 31192 19392 31195
rect 4989 31187 5190 31190
rect 615 31178 3797 31181
rect 615 31134 3750 31178
rect 3794 31134 3797 31178
rect 568 31131 3797 31134
rect 4989 31135 4992 31187
rect 5044 31135 5190 31187
rect 4989 31132 5190 31135
rect 14770 31187 14971 31190
rect 14770 31135 14916 31187
rect 14968 31135 14971 31187
rect 19342 31181 19345 31192
rect 14770 31132 14971 31135
rect 16163 31178 19345 31181
rect 16163 31134 16166 31178
rect 16210 31134 19345 31178
rect 19389 31134 19392 31192
rect 16163 31131 19392 31134
rect 5031 31096 5242 31099
rect 5031 31038 5034 31096
rect 5060 31038 5213 31096
rect 5239 31038 5242 31096
rect 5031 31035 5242 31038
rect 14718 31096 14929 31099
rect 14718 31038 14721 31096
rect 14747 31038 14900 31096
rect 14926 31038 14929 31096
rect 14718 31035 14929 31038
rect 504 30856 554 30859
rect 504 30798 507 30856
rect 551 30845 554 30856
rect 19406 30856 19456 30859
rect 19406 30845 19409 30856
rect 551 30842 3797 30845
rect 551 30798 3750 30842
rect 3794 30798 3797 30842
rect 504 30795 3797 30798
rect 16163 30842 19409 30845
rect 16163 30798 16166 30842
rect 16210 30798 19409 30842
rect 19453 30798 19456 30856
rect 16163 30795 19456 30798
rect 440 30792 490 30795
rect 440 30734 443 30792
rect 487 30781 490 30792
rect 19470 30792 19520 30795
rect 4989 30787 5190 30790
rect 487 30778 3797 30781
rect 487 30734 3750 30778
rect 3794 30734 3797 30778
rect 440 30731 3797 30734
rect 4989 30735 4992 30787
rect 5044 30735 5190 30787
rect 4989 30732 5190 30735
rect 14770 30787 14971 30790
rect 14770 30735 14916 30787
rect 14968 30735 14971 30787
rect 19470 30781 19473 30792
rect 14770 30732 14971 30735
rect 16163 30778 19473 30781
rect 16163 30734 16166 30778
rect 16210 30734 19473 30778
rect 19517 30734 19520 30792
rect 16163 30731 19520 30734
rect 5031 30696 5242 30699
rect 376 30655 426 30658
rect 376 30597 379 30655
rect 423 30644 426 30655
rect 423 30597 3588 30644
rect 5031 30638 5034 30696
rect 5060 30638 5213 30696
rect 5239 30638 5242 30696
rect 5031 30635 5242 30638
rect 14718 30696 14929 30699
rect 14718 30638 14721 30696
rect 14747 30638 14900 30696
rect 14926 30638 14929 30696
rect 19534 30655 19584 30658
rect 19534 30644 19537 30655
rect 14718 30635 14929 30638
rect 376 30594 3588 30597
rect 312 30591 362 30594
rect 312 30533 315 30591
rect 359 30580 362 30591
rect 359 30533 3518 30580
rect 312 30530 3518 30533
rect 40 30507 2858 30510
rect 40 30460 2811 30507
rect 2808 30449 2811 30460
rect 2855 30449 2858 30507
rect 2808 30446 2858 30449
rect 40 30417 2794 30420
rect 40 30370 2747 30417
rect 2744 30359 2747 30370
rect 2791 30359 2794 30417
rect 2744 30356 2794 30359
rect 3468 30381 3518 30530
rect 3538 30445 3588 30594
rect 5138 30618 5349 30621
rect 5138 30560 5141 30618
rect 5167 30560 5320 30618
rect 5346 30560 5349 30618
rect 5138 30557 5349 30560
rect 14611 30618 14822 30621
rect 14611 30560 14614 30618
rect 14640 30560 14793 30618
rect 14819 30560 14822 30618
rect 14611 30557 14822 30560
rect 16372 30597 19537 30644
rect 19581 30597 19584 30655
rect 16372 30594 19584 30597
rect 16372 30445 16422 30594
rect 19598 30591 19648 30594
rect 19598 30580 19601 30591
rect 3538 30442 3797 30445
rect 3538 30398 3750 30442
rect 3794 30398 3797 30442
rect 3538 30395 3797 30398
rect 16163 30442 16422 30445
rect 16163 30398 16166 30442
rect 16210 30398 16422 30442
rect 16163 30395 16422 30398
rect 16442 30533 19601 30580
rect 19645 30533 19648 30591
rect 16442 30530 19648 30533
rect 4989 30387 5190 30390
rect 3468 30378 3797 30381
rect 3468 30334 3750 30378
rect 3794 30334 3797 30378
rect 3468 30331 3797 30334
rect 4989 30335 4992 30387
rect 5044 30335 5190 30387
rect 4989 30332 5190 30335
rect 14770 30387 14971 30390
rect 14770 30335 14916 30387
rect 14968 30335 14971 30387
rect 16442 30381 16492 30530
rect 17102 30507 19920 30510
rect 17102 30449 17105 30507
rect 17149 30460 19920 30507
rect 17149 30449 17152 30460
rect 17102 30446 17152 30449
rect 14770 30332 14971 30335
rect 16163 30378 16492 30381
rect 16163 30334 16166 30378
rect 16210 30334 16492 30378
rect 17166 30417 19920 30420
rect 17166 30359 17169 30417
rect 17213 30370 19920 30417
rect 17213 30359 17216 30370
rect 17166 30356 17216 30359
rect 16163 30331 16492 30334
rect 5031 30296 5242 30299
rect 5031 30238 5034 30296
rect 5060 30238 5213 30296
rect 5239 30238 5242 30296
rect 5031 30235 5242 30238
rect 14718 30296 14929 30299
rect 14718 30238 14721 30296
rect 14747 30238 14900 30296
rect 14926 30238 14929 30296
rect 14718 30235 14929 30238
rect 248 30056 298 30059
rect 248 29998 251 30056
rect 295 30045 298 30056
rect 19662 30056 19712 30059
rect 19662 30045 19665 30056
rect 295 30042 3797 30045
rect 295 29998 3750 30042
rect 3794 29998 3797 30042
rect 248 29995 3797 29998
rect 16163 30042 19665 30045
rect 16163 29998 16166 30042
rect 16210 29998 19665 30042
rect 19709 29998 19712 30056
rect 16163 29995 19712 29998
rect 184 29992 234 29995
rect 184 29934 187 29992
rect 231 29981 234 29992
rect 19726 29992 19776 29995
rect 4989 29987 5190 29990
rect 231 29978 3797 29981
rect 231 29934 3750 29978
rect 3794 29934 3797 29978
rect 184 29931 3797 29934
rect 4989 29935 4992 29987
rect 5044 29935 5190 29987
rect 4989 29932 5190 29935
rect 14770 29987 14971 29990
rect 14770 29935 14916 29987
rect 14968 29935 14971 29987
rect 19726 29981 19729 29992
rect 14770 29932 14971 29935
rect 16163 29978 19729 29981
rect 16163 29934 16166 29978
rect 16210 29934 19729 29978
rect 19773 29934 19776 29992
rect 16163 29931 19776 29934
rect 5031 29896 5242 29899
rect 5031 29838 5034 29896
rect 5060 29838 5213 29896
rect 5239 29838 5242 29896
rect 5031 29835 5242 29838
rect 14718 29896 14929 29899
rect 14718 29838 14721 29896
rect 14747 29838 14900 29896
rect 14926 29838 14929 29896
rect 14718 29835 14929 29838
rect 5138 29818 5349 29821
rect 5138 29760 5141 29818
rect 5167 29760 5320 29818
rect 5346 29760 5349 29818
rect 5138 29757 5349 29760
rect 14611 29818 14822 29821
rect 14611 29760 14614 29818
rect 14640 29760 14793 29818
rect 14819 29760 14822 29818
rect 14611 29757 14822 29760
rect 3747 29642 3797 29645
rect 3747 29598 3750 29642
rect 3794 29598 3797 29642
rect 3747 29595 3797 29598
rect 16163 29642 16213 29645
rect 16163 29598 16166 29642
rect 16210 29598 16213 29642
rect 16163 29595 16213 29598
rect 4989 29587 5190 29590
rect 3747 29578 3797 29581
rect 3747 29534 3750 29578
rect 3794 29534 3797 29578
rect 3747 29531 3797 29534
rect 4989 29535 4992 29587
rect 5044 29535 5190 29587
rect 4989 29532 5190 29535
rect 14770 29587 14971 29590
rect 14770 29535 14916 29587
rect 14968 29535 14971 29587
rect 14770 29532 14971 29535
rect 16163 29578 16213 29581
rect 16163 29534 16166 29578
rect 16210 29534 16213 29578
rect 16163 29531 16213 29534
rect 5031 29496 5242 29499
rect 5031 29438 5034 29496
rect 5060 29438 5213 29496
rect 5239 29438 5242 29496
rect 5031 29435 5242 29438
rect 14718 29496 14929 29499
rect 14718 29438 14721 29496
rect 14747 29438 14900 29496
rect 14926 29438 14929 29496
rect 14718 29435 14929 29438
rect 3747 29242 3797 29245
rect 3747 29198 3750 29242
rect 3794 29198 3797 29242
rect 3747 29195 3797 29198
rect 16163 29242 16213 29245
rect 16163 29198 16166 29242
rect 16210 29198 16213 29242
rect 16163 29195 16213 29198
rect 4989 29187 5190 29190
rect 3747 29178 3797 29181
rect 3747 29134 3750 29178
rect 3794 29134 3797 29178
rect 3747 29131 3797 29134
rect 4989 29135 4992 29187
rect 5044 29135 5190 29187
rect 4989 29132 5190 29135
rect 14770 29187 14971 29190
rect 14770 29135 14916 29187
rect 14968 29135 14971 29187
rect 14770 29132 14971 29135
rect 16163 29178 16213 29181
rect 16163 29134 16166 29178
rect 16210 29134 16213 29178
rect 16163 29131 16213 29134
rect 5031 29096 5242 29099
rect 5031 29038 5034 29096
rect 5060 29038 5213 29096
rect 5239 29038 5242 29096
rect 5031 29035 5242 29038
rect 14718 29096 14929 29099
rect 14718 29038 14721 29096
rect 14747 29038 14900 29096
rect 14926 29038 14929 29096
rect 14718 29035 14929 29038
rect 40 29007 2730 29010
rect 40 28960 2683 29007
rect 2680 28949 2683 28960
rect 2727 28949 2730 29007
rect 17230 29007 19920 29010
rect 2680 28946 2730 28949
rect 5170 28997 5820 29000
rect 40 28917 2666 28920
rect 40 28870 2619 28917
rect 2616 28859 2619 28870
rect 2663 28859 2666 28917
rect 5170 28908 5175 28997
rect 5815 28908 5820 28997
rect 5170 28903 5820 28908
rect 14140 28998 14790 29003
rect 14140 28908 14145 28998
rect 14785 28908 14790 28998
rect 17230 28949 17233 29007
rect 17277 28960 19920 29007
rect 17277 28949 17280 28960
rect 17230 28946 17280 28949
rect 14140 28903 14790 28908
rect 17294 28917 19920 28920
rect 2616 28856 2666 28859
rect 17294 28859 17297 28917
rect 17341 28870 19920 28917
rect 17341 28859 17344 28870
rect 17294 28856 17344 28859
rect 40 27507 2602 27510
rect 40 27460 2555 27507
rect 2552 27449 2555 27460
rect 2599 27449 2602 27507
rect 2552 27446 2602 27449
rect 17358 27507 19920 27510
rect 17358 27449 17361 27507
rect 17405 27460 19920 27507
rect 17405 27449 17408 27460
rect 17358 27446 17408 27449
rect 40 27417 2538 27420
rect 40 27370 2491 27417
rect 2488 27359 2491 27370
rect 2535 27359 2538 27417
rect 2488 27356 2538 27359
rect 17422 27417 19920 27420
rect 17422 27359 17425 27417
rect 17469 27370 19920 27417
rect 17469 27359 17472 27370
rect 17422 27356 17472 27359
rect 40 26007 2474 26010
rect 40 25960 2427 26007
rect 2424 25949 2427 25960
rect 2471 25949 2474 26007
rect 2424 25946 2474 25949
rect 17486 26007 19920 26010
rect 17486 25949 17489 26007
rect 17533 25960 19920 26007
rect 17533 25949 17536 25960
rect 17486 25946 17536 25949
rect 40 25917 2410 25920
rect 40 25870 2363 25917
rect 2360 25859 2363 25870
rect 2407 25859 2410 25917
rect 2360 25856 2410 25859
rect 17550 25917 19920 25920
rect 17550 25859 17553 25917
rect 17597 25870 19920 25917
rect 17597 25859 17600 25870
rect 17550 25856 17600 25859
rect 40 24507 2346 24510
rect 40 24460 2299 24507
rect 2296 24449 2299 24460
rect 2343 24449 2346 24507
rect 2296 24446 2346 24449
rect 17614 24507 19920 24510
rect 17614 24449 17617 24507
rect 17661 24460 19920 24507
rect 17661 24449 17664 24460
rect 17614 24446 17664 24449
rect 40 24417 2282 24420
rect 40 24370 2235 24417
rect 2232 24359 2235 24370
rect 2279 24359 2282 24417
rect 2232 24356 2282 24359
rect 17678 24417 19920 24420
rect 17678 24359 17681 24417
rect 17725 24370 19920 24417
rect 17725 24359 17728 24370
rect 17678 24356 17728 24359
rect 40 23007 2218 23010
rect 40 22960 2171 23007
rect 2168 22949 2171 22960
rect 2215 22949 2218 23007
rect 2168 22946 2218 22949
rect 17742 23007 19920 23010
rect 17742 22949 17745 23007
rect 17789 22960 19920 23007
rect 17789 22949 17792 22960
rect 17742 22946 17792 22949
rect 40 22917 2154 22920
rect 40 22870 2107 22917
rect 2104 22859 2107 22870
rect 2151 22859 2154 22917
rect 2104 22856 2154 22859
rect 17806 22917 19920 22920
rect 17806 22859 17809 22917
rect 17853 22870 19920 22917
rect 17853 22859 17856 22870
rect 17806 22856 17856 22859
rect 40 21507 2090 21510
rect 40 21460 2043 21507
rect 2040 21449 2043 21460
rect 2087 21449 2090 21507
rect 2040 21446 2090 21449
rect 17870 21507 19920 21510
rect 17870 21449 17873 21507
rect 17917 21460 19920 21507
rect 17917 21449 17920 21460
rect 17870 21446 17920 21449
rect 40 21417 2026 21420
rect 40 21370 1979 21417
rect 1976 21359 1979 21370
rect 2023 21359 2026 21417
rect 1976 21356 2026 21359
rect 17934 21417 19920 21420
rect 17934 21359 17937 21417
rect 17981 21370 19920 21417
rect 17981 21359 17984 21370
rect 17934 21356 17984 21359
rect 40 20007 1962 20010
rect 40 19960 1915 20007
rect 1912 19949 1915 19960
rect 1959 19949 1962 20007
rect 1912 19946 1962 19949
rect 17998 20007 19920 20010
rect 17998 19949 18001 20007
rect 18045 19960 19920 20007
rect 18045 19949 18048 19960
rect 17998 19946 18048 19949
rect 40 19917 1898 19920
rect 40 19870 1851 19917
rect 1848 19859 1851 19870
rect 1895 19859 1898 19917
rect 1848 19856 1898 19859
rect 18062 19917 19920 19920
rect 18062 19859 18065 19917
rect 18109 19870 19920 19917
rect 18109 19859 18112 19870
rect 18062 19856 18112 19859
rect 40 18507 1834 18510
rect 40 18460 1787 18507
rect 1784 18449 1787 18460
rect 1831 18449 1834 18507
rect 1784 18446 1834 18449
rect 18126 18507 19920 18510
rect 18126 18449 18129 18507
rect 18173 18460 19920 18507
rect 18173 18449 18176 18460
rect 18126 18446 18176 18449
rect 40 18417 1770 18420
rect 40 18370 1723 18417
rect 1720 18359 1723 18370
rect 1767 18359 1770 18417
rect 1720 18356 1770 18359
rect 18190 18417 19920 18420
rect 18190 18359 18193 18417
rect 18237 18370 19920 18417
rect 18237 18359 18240 18370
rect 18190 18356 18240 18359
rect 40 17007 1706 17010
rect 40 16960 1659 17007
rect 1656 16949 1659 16960
rect 1703 16949 1706 17007
rect 1656 16946 1706 16949
rect 18254 17007 19920 17010
rect 18254 16949 18257 17007
rect 18301 16960 19920 17007
rect 18301 16949 18304 16960
rect 18254 16946 18304 16949
rect 40 16917 1642 16920
rect 40 16870 1595 16917
rect 1592 16859 1595 16870
rect 1639 16859 1642 16917
rect 1592 16856 1642 16859
rect 18318 16917 19920 16920
rect 18318 16859 18321 16917
rect 18365 16870 19920 16917
rect 18365 16859 18368 16870
rect 18318 16856 18368 16859
rect 40 15507 1578 15510
rect 40 15460 1531 15507
rect 1528 15449 1531 15460
rect 1575 15449 1578 15507
rect 1528 15446 1578 15449
rect 18382 15507 19920 15510
rect 18382 15449 18385 15507
rect 18429 15460 19920 15507
rect 18429 15449 18432 15460
rect 18382 15446 18432 15449
rect 40 15417 1514 15420
rect 40 15370 1467 15417
rect 1464 15359 1467 15370
rect 1511 15359 1514 15417
rect 1464 15356 1514 15359
rect 18446 15417 19920 15420
rect 18446 15359 18449 15417
rect 18493 15370 19920 15417
rect 18493 15359 18496 15370
rect 18446 15356 18496 15359
rect 40 14007 1450 14010
rect 40 13960 1403 14007
rect 1400 13949 1403 13960
rect 1447 13949 1450 14007
rect 1400 13946 1450 13949
rect 18510 14007 19920 14010
rect 18510 13949 18513 14007
rect 18557 13960 19920 14007
rect 18557 13949 18560 13960
rect 18510 13946 18560 13949
rect 40 13917 1386 13920
rect 40 13870 1339 13917
rect 1336 13859 1339 13870
rect 1383 13859 1386 13917
rect 1336 13856 1386 13859
rect 18574 13917 19920 13920
rect 18574 13859 18577 13917
rect 18621 13870 19920 13917
rect 18621 13859 18624 13870
rect 18574 13856 18624 13859
rect 40 12507 1322 12510
rect 40 12460 1275 12507
rect 1272 12449 1275 12460
rect 1319 12449 1322 12507
rect 1272 12446 1322 12449
rect 18638 12507 19920 12510
rect 18638 12449 18641 12507
rect 18685 12460 19920 12507
rect 18685 12449 18688 12460
rect 18638 12446 18688 12449
rect 40 12417 1258 12420
rect 40 12370 1211 12417
rect 1208 12359 1211 12370
rect 1255 12359 1258 12417
rect 1208 12356 1258 12359
rect 18702 12417 19920 12420
rect 18702 12359 18705 12417
rect 18749 12370 19920 12417
rect 18749 12359 18752 12370
rect 18702 12356 18752 12359
rect 40 11007 1194 11010
rect 40 10960 1147 11007
rect 1144 10949 1147 10960
rect 1191 10949 1194 11007
rect 1144 10946 1194 10949
rect 18766 11007 19920 11010
rect 18766 10949 18769 11007
rect 18813 10960 19920 11007
rect 18813 10949 18816 10960
rect 18766 10946 18816 10949
rect 40 10917 1130 10920
rect 40 10870 1083 10917
rect 1080 10859 1083 10870
rect 1127 10859 1130 10917
rect 1080 10856 1130 10859
rect 18830 10917 19920 10920
rect 18830 10859 18833 10917
rect 18877 10870 19920 10917
rect 18877 10859 18880 10870
rect 18830 10856 18880 10859
rect 40 9507 1066 9510
rect 40 9460 1019 9507
rect 1016 9449 1019 9460
rect 1063 9449 1066 9507
rect 1016 9446 1066 9449
rect 18894 9507 19920 9510
rect 18894 9449 18897 9507
rect 18941 9460 19920 9507
rect 18941 9449 18944 9460
rect 18894 9446 18944 9449
rect 40 9417 1002 9420
rect 40 9370 955 9417
rect 952 9359 955 9370
rect 999 9359 1002 9417
rect 952 9356 1002 9359
rect 18958 9417 19920 9420
rect 18958 9359 18961 9417
rect 19005 9370 19920 9417
rect 19005 9359 19008 9370
rect 18958 9356 19008 9359
rect 40 8007 938 8010
rect 40 7960 891 8007
rect 888 7949 891 7960
rect 935 7949 938 8007
rect 888 7946 938 7949
rect 19022 8007 19920 8010
rect 19022 7949 19025 8007
rect 19069 7960 19920 8007
rect 19069 7949 19072 7960
rect 19022 7946 19072 7949
rect 40 7917 874 7920
rect 40 7870 827 7917
rect 824 7859 827 7870
rect 871 7859 874 7917
rect 824 7856 874 7859
rect 19086 7917 19920 7920
rect 19086 7859 19089 7917
rect 19133 7870 19920 7917
rect 19133 7859 19136 7870
rect 19086 7856 19136 7859
rect 40 6507 810 6510
rect 40 6460 763 6507
rect 760 6449 763 6460
rect 807 6449 810 6507
rect 760 6446 810 6449
rect 19150 6507 19920 6510
rect 19150 6449 19153 6507
rect 19197 6460 19920 6507
rect 19197 6449 19200 6460
rect 19150 6446 19200 6449
rect 40 6417 746 6420
rect 40 6370 699 6417
rect 696 6359 699 6370
rect 743 6359 746 6417
rect 696 6356 746 6359
rect 19214 6417 19920 6420
rect 19214 6359 19217 6417
rect 19261 6370 19920 6417
rect 19261 6359 19264 6370
rect 19214 6356 19264 6359
rect 8774 6201 12968 6204
rect 8774 6199 12871 6201
rect 8774 6109 8779 6199
rect 8969 6109 12871 6199
rect 8774 6107 12871 6109
rect 12965 6107 12968 6201
rect 8774 6104 12968 6107
rect 9042 6033 13106 6036
rect 9042 6031 13009 6033
rect 9042 5941 9047 6031
rect 9237 5941 13009 6031
rect 9042 5939 13009 5941
rect 13103 5939 13106 6033
rect 9042 5936 13106 5939
rect 9310 5865 13244 5868
rect 9310 5863 13147 5865
rect 9310 5773 9315 5863
rect 9505 5773 13147 5863
rect 9310 5771 13147 5773
rect 13241 5771 13244 5865
rect 9310 5768 13244 5771
rect 9578 5697 13382 5700
rect 9578 5695 13285 5697
rect 9578 5605 9583 5695
rect 9773 5605 13285 5695
rect 9578 5603 13285 5605
rect 13379 5603 13382 5697
rect 9578 5600 13382 5603
rect 12868 5577 12968 5580
rect 12868 5483 12871 5577
rect 12965 5483 12968 5577
rect 12868 5480 12968 5483
rect 13006 5577 13106 5580
rect 13006 5483 13009 5577
rect 13103 5483 13106 5577
rect 13006 5480 13106 5483
rect 13144 5577 13244 5580
rect 13144 5483 13147 5577
rect 13241 5483 13244 5577
rect 13144 5480 13244 5483
rect 40 5007 682 5010
rect 40 4960 635 5007
rect 632 4949 635 4960
rect 679 4949 682 5007
rect 632 4946 682 4949
rect 19278 5007 19920 5010
rect 19278 4949 19281 5007
rect 19325 4960 19920 5007
rect 19325 4949 19328 4960
rect 19278 4946 19328 4949
rect 40 4917 618 4920
rect 40 4870 571 4917
rect 568 4859 571 4870
rect 615 4859 618 4917
rect 568 4856 618 4859
rect 19342 4917 19920 4920
rect 19342 4859 19345 4917
rect 19389 4870 19920 4917
rect 19389 4859 19392 4870
rect 19342 4856 19392 4859
rect 40 3507 554 3510
rect 40 3460 507 3507
rect 504 3449 507 3460
rect 551 3449 554 3507
rect 504 3446 554 3449
rect 19406 3507 19920 3510
rect 19406 3449 19409 3507
rect 19453 3460 19920 3507
rect 19453 3449 19456 3460
rect 19406 3446 19456 3449
rect 40 3417 490 3420
rect 40 3370 443 3417
rect 440 3359 443 3370
rect 487 3359 490 3417
rect 440 3356 490 3359
rect 19470 3417 19920 3420
rect 19470 3359 19473 3417
rect 19517 3370 19920 3417
rect 19517 3359 19520 3370
rect 19470 3356 19520 3359
rect 6811 2156 6869 2159
rect 6811 2130 6814 2156
rect 6866 2130 6869 2156
rect 6083 2049 6141 2052
rect 6083 2023 6086 2049
rect 6138 2023 6141 2049
rect 40 2007 426 2010
rect 40 1960 379 2007
rect 376 1949 379 1960
rect 423 1949 426 2007
rect 376 1946 426 1949
rect 40 1917 362 1920
rect 40 1870 315 1917
rect 312 1859 315 1870
rect 359 1859 362 1917
rect 312 1856 362 1859
rect 6083 1870 6141 2023
rect 6083 1844 6086 1870
rect 6138 1844 6141 1870
rect 6083 1841 6141 1844
rect 6483 2049 6541 2052
rect 6483 2023 6486 2049
rect 6538 2023 6541 2049
rect 6483 1870 6541 2023
rect 6811 1977 6869 2130
rect 7611 2156 7669 2159
rect 7611 2130 7614 2156
rect 7666 2130 7669 2156
rect 6811 1951 6814 1977
rect 6866 1951 6869 1977
rect 6811 1948 6869 1951
rect 6883 2049 6941 2052
rect 6883 2023 6886 2049
rect 6938 2023 6941 2049
rect 6483 1844 6486 1870
rect 6538 1844 6541 1870
rect 6483 1841 6541 1844
rect 6883 1870 6941 2023
rect 6883 1844 6886 1870
rect 6938 1844 6941 1870
rect 6883 1841 6941 1844
rect 7283 2049 7341 2052
rect 7283 2023 7286 2049
rect 7338 2023 7341 2049
rect 7283 1870 7341 2023
rect 7611 1977 7669 2130
rect 8411 2156 8469 2159
rect 8411 2130 8414 2156
rect 8466 2130 8469 2156
rect 7611 1951 7614 1977
rect 7666 1951 7669 1977
rect 7611 1948 7669 1951
rect 7683 2049 7741 2052
rect 7683 2023 7686 2049
rect 7738 2023 7741 2049
rect 7283 1844 7286 1870
rect 7338 1844 7341 1870
rect 7283 1841 7341 1844
rect 7683 1870 7741 2023
rect 7683 1844 7686 1870
rect 7738 1844 7741 1870
rect 7683 1841 7741 1844
rect 8083 2049 8141 2052
rect 8083 2023 8086 2049
rect 8138 2023 8141 2049
rect 8083 1870 8141 2023
rect 8411 1977 8469 2130
rect 9211 2156 9269 2159
rect 9211 2130 9214 2156
rect 9266 2130 9269 2156
rect 8411 1951 8414 1977
rect 8466 1951 8469 1977
rect 8411 1948 8469 1951
rect 8483 2049 8541 2052
rect 8483 2023 8486 2049
rect 8538 2023 8541 2049
rect 8083 1844 8086 1870
rect 8138 1844 8141 1870
rect 8083 1841 8141 1844
rect 8483 1870 8541 2023
rect 8483 1844 8486 1870
rect 8538 1844 8541 1870
rect 8483 1841 8541 1844
rect 8883 2049 8941 2052
rect 8883 2023 8886 2049
rect 8938 2023 8941 2049
rect 8883 1870 8941 2023
rect 9211 1977 9269 2130
rect 10011 2156 10069 2159
rect 10011 2130 10014 2156
rect 10066 2130 10069 2156
rect 9211 1951 9214 1977
rect 9266 1951 9269 1977
rect 9211 1948 9269 1951
rect 9283 2049 9341 2052
rect 9283 2023 9286 2049
rect 9338 2023 9341 2049
rect 8883 1844 8886 1870
rect 8938 1844 8941 1870
rect 8883 1841 8941 1844
rect 9283 1870 9341 2023
rect 9283 1844 9286 1870
rect 9338 1844 9341 1870
rect 9283 1841 9341 1844
rect 9683 2049 9741 2052
rect 9683 2023 9686 2049
rect 9738 2023 9741 2049
rect 9683 1870 9741 2023
rect 10011 1977 10069 2130
rect 10811 2156 10869 2159
rect 10811 2130 10814 2156
rect 10866 2130 10869 2156
rect 10011 1951 10014 1977
rect 10066 1951 10069 1977
rect 10011 1948 10069 1951
rect 10083 2049 10141 2052
rect 10083 2023 10086 2049
rect 10138 2023 10141 2049
rect 9683 1844 9686 1870
rect 9738 1844 9741 1870
rect 9683 1841 9741 1844
rect 10083 1870 10141 2023
rect 10083 1844 10086 1870
rect 10138 1844 10141 1870
rect 10083 1841 10141 1844
rect 10483 2049 10541 2052
rect 10483 2023 10486 2049
rect 10538 2023 10541 2049
rect 10483 1870 10541 2023
rect 10811 1977 10869 2130
rect 11611 2156 11669 2159
rect 11611 2130 11614 2156
rect 11666 2130 11669 2156
rect 10811 1951 10814 1977
rect 10866 1951 10869 1977
rect 10811 1948 10869 1951
rect 10883 2049 10941 2052
rect 10883 2023 10886 2049
rect 10938 2023 10941 2049
rect 10483 1844 10486 1870
rect 10538 1844 10541 1870
rect 10483 1841 10541 1844
rect 10883 1870 10941 2023
rect 10883 1844 10886 1870
rect 10938 1844 10941 1870
rect 10883 1841 10941 1844
rect 11283 2049 11341 2052
rect 11283 2023 11286 2049
rect 11338 2023 11341 2049
rect 11283 1870 11341 2023
rect 11611 1977 11669 2130
rect 11611 1951 11614 1977
rect 11666 1951 11669 1977
rect 11611 1948 11669 1951
rect 11683 2049 11741 2052
rect 11683 2023 11686 2049
rect 11738 2023 11741 2049
rect 11283 1844 11286 1870
rect 11338 1844 11341 1870
rect 11283 1841 11341 1844
rect 11683 1870 11741 2023
rect 11683 1844 11686 1870
rect 11738 1844 11741 1870
rect 11683 1841 11741 1844
rect 12083 2049 12141 2052
rect 12083 2023 12086 2049
rect 12138 2023 12141 2049
rect 12083 1870 12141 2023
rect 12440 1977 12520 2130
rect 12440 1903 12443 1977
rect 12517 1903 12520 1977
rect 19534 2007 19920 2010
rect 19534 1949 19537 2007
rect 19581 1960 19920 2007
rect 19581 1949 19584 1960
rect 19534 1946 19584 1949
rect 12440 1900 12520 1903
rect 19598 1917 19920 1920
rect 12083 1844 12086 1870
rect 12138 1844 12141 1870
rect 19598 1859 19601 1917
rect 19645 1870 19920 1917
rect 19645 1859 19648 1870
rect 19598 1856 19648 1859
rect 12083 1841 12141 1844
rect 40 507 298 510
rect 40 460 251 507
rect 248 449 251 460
rect 295 449 298 507
rect 248 446 298 449
rect 19662 507 19920 510
rect 19662 449 19665 507
rect 19709 460 19920 507
rect 19709 449 19712 460
rect 19662 446 19712 449
rect 40 417 234 420
rect 40 370 187 417
rect 184 359 187 370
rect 231 359 234 417
rect 184 356 234 359
rect 19726 417 19920 420
rect 19726 359 19729 417
rect 19773 370 19920 417
rect 19773 359 19776 370
rect 19726 356 19776 359
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -220 -5 -140 0
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect -220 -80 -140 -75
rect 20100 -5 20180 0
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
rect -14 -110 19973 -107
rect -14 -136 -11 -110
rect 15 -136 12250 -110
rect 12276 -136 19944 -110
rect 19970 -136 19973 -110
rect -14 -139 19973 -136
rect -268 -156 20227 -153
rect -268 -182 -265 -156
rect -239 -182 12196 -156
rect 12222 -182 20198 -156
rect 20224 -182 20227 -156
rect -268 -185 20227 -182
rect -2016 -202 21975 -199
rect -2016 -228 -2011 -202
rect -1985 -228 11850 -202
rect 11876 -228 21944 -202
rect 21970 -228 21975 -202
rect -2016 -231 21975 -228
rect -2270 -248 22229 -245
rect -2270 -274 -2265 -248
rect -2239 -274 11796 -248
rect 11822 -274 22198 -248
rect 22224 -274 22229 -248
rect -2270 -277 22229 -274
rect -4016 -294 23975 -291
rect -4016 -320 -4011 -294
rect -3985 -320 11450 -294
rect 11476 -320 23944 -294
rect 23970 -320 23975 -294
rect -4016 -323 23975 -320
rect -4270 -340 24229 -337
rect -4270 -366 -4265 -340
rect -4239 -366 11396 -340
rect 11422 -366 24198 -340
rect 24224 -366 24229 -340
rect -4270 -369 24229 -366
rect -6016 -386 25975 -383
rect -6016 -412 -6011 -386
rect -5985 -412 11050 -386
rect 11076 -412 25944 -386
rect 25970 -412 25975 -386
rect -6016 -415 25975 -412
rect -6270 -432 26229 -429
rect -6270 -458 -6265 -432
rect -6239 -458 10996 -432
rect 11022 -458 26198 -432
rect 26224 -458 26229 -432
rect -6270 -461 26229 -458
rect -8016 -478 27975 -475
rect -8016 -504 -8011 -478
rect -7985 -504 10650 -478
rect 10676 -504 27944 -478
rect 27970 -504 27975 -478
rect -8016 -507 27975 -504
rect -8270 -524 28229 -521
rect -8270 -550 -8265 -524
rect -8239 -550 10596 -524
rect 10622 -550 28198 -524
rect 28224 -550 28229 -524
rect -8270 -553 28229 -550
rect -10016 -570 29975 -567
rect -10016 -596 -10011 -570
rect -9985 -596 10250 -570
rect 10276 -596 29944 -570
rect 29970 -596 29975 -570
rect -10016 -599 29975 -596
rect -10270 -616 30229 -613
rect -10270 -642 -10265 -616
rect -10239 -642 10196 -616
rect 10222 -642 30198 -616
rect 30224 -642 30229 -616
rect -10270 -645 30229 -642
rect -12016 -662 31975 -659
rect -12016 -688 -12011 -662
rect -11985 -688 9850 -662
rect 9876 -688 31944 -662
rect 31970 -688 31975 -662
rect -12016 -691 31975 -688
rect -12270 -708 32229 -705
rect -12270 -734 -12265 -708
rect -12239 -734 9796 -708
rect 9822 -734 32198 -708
rect 32224 -734 32229 -708
rect -12270 -737 32229 -734
rect -14016 -754 33975 -751
rect -14016 -780 -14011 -754
rect -13985 -780 9450 -754
rect 9476 -780 33944 -754
rect 33970 -780 33975 -754
rect -14016 -783 33975 -780
rect -14270 -800 34229 -797
rect -14270 -826 -14265 -800
rect -14239 -826 9396 -800
rect 9422 -826 34198 -800
rect 34224 -826 34229 -800
rect -14270 -829 34229 -826
rect -16014 -846 35973 -843
rect -16014 -872 -16011 -846
rect -15985 -872 9050 -846
rect 9076 -872 35944 -846
rect 35970 -872 35973 -846
rect -16014 -875 35973 -872
rect -16268 -892 36227 -889
rect -16268 -918 -16265 -892
rect -16239 -918 8996 -892
rect 9022 -918 36198 -892
rect 36224 -918 36227 -892
rect -16268 -921 36227 -918
rect -18014 -938 37973 -935
rect -18014 -964 -18011 -938
rect -17985 -964 8650 -938
rect 8676 -964 37944 -938
rect 37970 -964 37973 -938
rect -18014 -967 37973 -964
rect -18268 -984 38229 -981
rect -18268 -1010 -18265 -984
rect -18239 -1010 8596 -984
rect 8622 -1010 38198 -984
rect 38224 -1010 38229 -984
rect -18268 -1013 38229 -1010
<< via2 >>
rect 10923 42777 11113 42867
rect 10655 42639 10845 42729
rect 10387 42501 10577 42591
rect 10119 42363 10309 42453
rect 9851 42225 10041 42315
rect 5325 41787 5815 41877
rect 14145 41787 14635 41877
rect 5175 28908 5815 28997
rect 14145 28997 14785 28998
rect 14145 28908 14785 28997
rect 8779 6109 8969 6199
rect 9047 5941 9237 6031
rect 9315 5773 9505 5863
rect 9583 5605 9773 5695
rect -18215 -75 -18145 -5
rect -16215 -75 -16145 -5
rect -14215 -75 -14145 -5
rect -12215 -75 -12145 -5
rect -10215 -75 -10145 -5
rect -8215 -75 -8145 -5
rect -6215 -75 -6145 -5
rect -4215 -75 -4145 -5
rect -2215 -75 -2145 -5
rect -215 -75 -145 -5
rect 20105 -75 20175 -5
rect 22105 -75 22175 -5
rect 24105 -75 24175 -5
rect 26105 -75 26175 -5
rect 28105 -75 28175 -5
rect 30105 -75 30175 -5
rect 32105 -75 32175 -5
rect 34105 -75 34175 -5
rect 36105 -75 36175 -5
rect 38105 -75 38175 -5
<< metal3 >>
rect 5100 44900 5900 45000
rect 6100 44800 6900 45000
rect 6100 44430 6130 44800
rect 6870 44430 6900 44800
rect 6100 44420 6900 44430
rect 7300 43600 7500 45000
rect 7900 43900 8100 45000
rect 8500 44200 8700 45000
rect 9100 44500 9300 45000
rect 9700 44800 9900 45000
rect 9700 44600 10046 44800
rect 10300 44620 10500 45000
rect 9100 44300 9778 44500
rect 8500 44000 9510 44200
rect 7900 43700 9242 43900
rect 7300 43400 8974 43600
rect 5320 41877 5820 41882
rect 5320 41787 5325 41877
rect 5815 41787 5820 41877
rect 5320 41782 5820 41787
rect 5170 28998 5820 29001
rect 5170 28908 5175 28998
rect 5815 28908 5820 28998
rect 5170 28903 5820 28908
rect 8774 6199 8974 43400
rect 8774 6109 8779 6199
rect 8969 6109 8974 6199
rect 8774 6104 8974 6109
rect 9042 6031 9242 43700
rect 9042 5941 9047 6031
rect 9237 5941 9242 6031
rect 9042 5936 9242 5941
rect 9310 5863 9510 44000
rect 9310 5773 9315 5863
rect 9505 5773 9510 5863
rect 9310 5768 9510 5773
rect 9578 5695 9778 44300
rect 9846 42315 10046 44600
rect 10114 44420 10500 44620
rect 10114 42453 10314 44420
rect 10900 44320 11100 45000
rect 10382 44120 11100 44320
rect 10382 42591 10582 44120
rect 11500 44020 11700 45000
rect 10650 43820 11700 44020
rect 10650 42729 10850 43820
rect 12100 43720 12300 45000
rect 12700 44900 13500 45000
rect 13700 44800 14500 45000
rect 13700 44430 13730 44800
rect 14470 44430 14500 44800
rect 13700 44420 14500 44430
rect 10918 43520 12300 43720
rect 10918 42867 11118 43520
rect 10918 42777 10923 42867
rect 11113 42777 11118 42867
rect 10918 42772 11118 42777
rect 10650 42639 10655 42729
rect 10845 42639 10850 42729
rect 10650 42634 10850 42639
rect 10382 42501 10387 42591
rect 10577 42501 10582 42591
rect 10382 42496 10582 42501
rect 10114 42363 10119 42453
rect 10309 42363 10314 42453
rect 10114 42358 10314 42363
rect 9846 42225 9851 42315
rect 10041 42225 10046 42315
rect 9846 42220 10046 42225
rect 14140 41877 14640 41882
rect 14140 41787 14145 41877
rect 14635 41787 14640 41877
rect 14140 41782 14640 41787
rect 14140 28998 14790 29003
rect 14140 28908 14145 28998
rect 14785 28908 14790 28998
rect 14140 28903 14790 28908
rect 9578 5605 9583 5695
rect 9773 5605 9778 5695
rect 9578 5600 9778 5605
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -220 -5 -140 0
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect -220 -80 -140 -75
rect 20100 -5 20180 0
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
<< via3 >>
rect 6130 44430 6870 44800
rect 5325 41787 5815 41877
rect 5175 28997 5815 28998
rect 5175 28908 5815 28997
rect 13730 44430 14470 44800
rect 14145 41787 14635 41877
rect 14145 28908 14785 28998
<< metal4 >>
rect 6100 44800 14500 44801
rect 5000 44430 6130 44800
rect 6870 44430 13730 44800
rect 14470 44430 14900 44800
rect 5000 44400 14900 44430
rect 5000 41877 6200 44400
rect 5000 41787 5325 41877
rect 5815 41787 6200 41877
rect 5000 28998 6200 41787
rect 5000 28908 5175 28998
rect 5815 28908 6200 28998
rect 5000 28900 6200 28908
rect 13700 41877 14900 44400
rect 13700 41787 14145 41877
rect 14635 41787 14900 41877
rect 13700 28998 14900 41787
rect 13700 28908 14145 28998
rect 14785 28908 14900 28998
rect 13700 28900 14900 28908
<< via4 >>
rect -18900 -380 -18300 -80
rect -16900 -380 -16300 -80
rect -14900 -380 -14300 -80
rect -12900 -380 -12300 -80
rect -10900 -380 -10300 -80
rect -8900 -380 -8300 -80
rect -6900 -380 -6300 -80
rect -4900 -380 -4300 -80
rect -2900 -380 -2300 -80
rect -900 -380 -300 -80
rect 20920 -380 21520 -80
rect 22920 -380 23520 -80
rect 24920 -380 25520 -80
rect 26920 -380 27520 -80
rect 28920 -380 29520 -80
rect 30920 -380 31520 -80
rect 32920 -380 33520 -80
rect 34920 -380 35520 -80
rect 36920 -380 37520 -80
rect 38920 -380 39520 -80
<< metal5 >>
rect -19900 -600 -19300 0
rect -18900 -60 -18300 0
rect -18920 -80 -18280 -60
rect -18920 -380 -18900 -80
rect -18300 -380 -18280 -80
rect -18920 -400 -18280 -380
rect -17900 -600 -17300 0
rect -16900 -60 -16300 0
rect -16920 -80 -16280 -60
rect -16920 -380 -16900 -80
rect -16300 -380 -16280 -80
rect -16920 -400 -16280 -380
rect -15900 -600 -15300 0
rect -14900 -60 -14300 0
rect -14920 -80 -14280 -60
rect -14920 -380 -14900 -80
rect -14300 -380 -14280 -80
rect -14920 -400 -14280 -380
rect -13900 -600 -13300 0
rect -12900 -60 -12300 0
rect -12920 -80 -12280 -60
rect -12920 -380 -12900 -80
rect -12300 -380 -12280 -80
rect -12920 -400 -12280 -380
rect -11900 -600 -11300 0
rect -10900 -60 -10300 0
rect -10920 -80 -10280 -60
rect -10920 -380 -10900 -80
rect -10300 -380 -10280 -80
rect -10920 -400 -10280 -380
rect -9900 -600 -9300 0
rect -8900 -60 -8300 0
rect -8920 -80 -8280 -60
rect -8920 -380 -8900 -80
rect -8300 -380 -8280 -80
rect -8920 -400 -8280 -380
rect -7900 -600 -7300 0
rect -6900 -60 -6300 0
rect -6920 -80 -6280 -60
rect -6920 -380 -6900 -80
rect -6300 -380 -6280 -80
rect -6920 -400 -6280 -380
rect -5900 -600 -5300 0
rect -4900 -60 -4300 0
rect -4920 -80 -4280 -60
rect -4920 -380 -4900 -80
rect -4300 -380 -4280 -80
rect -4920 -400 -4280 -380
rect -3900 -600 -3300 0
rect -2900 -60 -2300 0
rect -2920 -80 -2280 -60
rect -2920 -380 -2900 -80
rect -2300 -380 -2280 -80
rect -2920 -400 -2280 -380
rect -1900 -600 -1300 0
rect -900 -60 -300 0
rect -920 -80 -280 -60
rect -920 -380 -900 -80
rect -300 -380 -280 -80
rect -920 -400 -280 -380
rect 19920 -600 20520 0
rect 20920 -60 21520 0
rect 20900 -80 21540 -60
rect 20900 -380 20920 -80
rect 21520 -380 21540 -80
rect 20900 -400 21540 -380
rect 21920 -600 22520 0
rect 22920 -60 23520 0
rect 22900 -80 23540 -60
rect 22900 -380 22920 -80
rect 23520 -380 23540 -80
rect 22900 -400 23540 -380
rect 23920 -600 24520 0
rect 24920 -60 25520 0
rect 24900 -80 25540 -60
rect 24900 -380 24920 -80
rect 25520 -380 25540 -80
rect 24900 -400 25540 -380
rect 25920 -600 26520 0
rect 26920 -60 27520 0
rect 26900 -80 27540 -60
rect 26900 -380 26920 -80
rect 27520 -380 27540 -80
rect 26900 -400 27540 -380
rect 27920 -600 28520 0
rect 28920 -60 29520 0
rect 28900 -80 29540 -60
rect 28900 -380 28920 -80
rect 29520 -380 29540 -80
rect 28900 -400 29540 -380
rect 29920 -600 30520 0
rect 30920 -60 31520 0
rect 30900 -80 31540 -60
rect 30900 -380 30920 -80
rect 31520 -380 31540 -80
rect 30900 -400 31540 -380
rect 31920 -600 32520 0
rect 32920 -60 33520 0
rect 32900 -80 33540 -60
rect 32900 -380 32920 -80
rect 33520 -380 33540 -80
rect 32900 -400 33540 -380
rect 33920 -600 34520 0
rect 34920 -60 35520 0
rect 34900 -80 35540 -60
rect 34900 -380 34920 -80
rect 35520 -380 35540 -80
rect 34900 -400 35540 -380
rect 35920 -600 36520 0
rect 36920 -60 37520 0
rect 36900 -80 37540 -60
rect 36900 -380 36920 -80
rect 37520 -380 37540 -80
rect 36900 -400 37540 -380
rect 37920 -600 38520 0
rect 38920 -60 39520 0
rect 38900 -80 39540 -60
rect 38900 -380 38920 -80
rect 39520 -380 39540 -80
rect 38900 -400 39540 -380
rect -19900 -1400 38520 -600
use array_column_decode  array_column_decode_0
timestamp 1717473404
transform 0 1 -520 -1 0 3560
box -2020 6520 1560 13936
use array_core_block0  array_core_block0_0
timestamp 1717516356
transform 1 0 -20000 0 1 30696
box -33 -696 19983 14118
use array_core_block1  array_core_block1_0
timestamp 1717516447
transform 1 0 -20000 0 1 15000
box -33 0 19983 14814
use array_core_block2  array_core_block2_0
timestamp 1717516403
transform 1 0 -20000 0 1 0
box -33 0 19983 14819
use array_core_block3  array_core_block3_0
timestamp 1717473404
transform -1 0 39983 0 -1 44411
box -33 0 19983 14411
use array_core_block4  array_core_block4_0
timestamp 1717473404
transform -1 0 39983 0 -1 29411
box -33 0 19983 14411
use array_core_block5  array_core_block5_0
timestamp 1717473404
transform -1 0 39983 0 1 0
box -33 0 19983 14623
use array_core_block_mirrored_routing  array_core_block_mirrored_routing_0
array 0 0 19940 0 2 15000
timestamp 1717473404
transform 1 0 19020 0 1 0
box 900 0 20840 15000
use array_core_block_routing  array_core_block_routing_1
array 0 0 19760 0 2 15000
timestamp 1717473404
transform 1 0 -20800 0 1 0
box 800 0 20840 15000
use array_row_decode  array_row_decode_0
timestamp 1717473404
transform 1 0 13210 0 1 28832
box -2020 168 1560 14074
use array_row_decode  array_row_decode_1
timestamp 1717473404
transform -1 0 6750 0 1 28832
box -2020 168 1560 14074
use lsi1v8o5v0  lsi1v8o5v0_0
array 0 0 1161 0 31 -400
timestamp 1717473404
transform -1 0 5048 0 -1 29307
box -42 -60 1301 293
use lsi1v8o5v0  lsi1v8o5v0_1
array 0 0 1161 0 31 -400
timestamp 1717473404
transform 1 0 14912 0 -1 29307
box -42 -60 1301 293
use lsi1v8o5v0  lsi1v8o5v0_2
array 0 0 1161 0 15 -400
timestamp 1717473404
transform 0 -1 6355 -1 0 1858
box -42 -60 1301 293
use tg5v0  tg5v0_0
array 0 0 -800 0 9 2000
timestamp 1717473404
transform 0 -1 90 -1 0 -983
box 14 0 817 445
use tg5v0  tg5v0_1
array 0 0 -800 0 9 2000
timestamp 1717473404
transform 0 1 19869 -1 0 -983
box 14 0 817 445
<< labels >>
flabel metal3 7300 44900 7500 45000 0 FreeSans 400 0 0 0 a[0]
port 3 nsew
flabel metal3 7900 44900 8100 45000 0 FreeSans 400 0 0 0 a[1]
port 4 nsew signal input
flabel metal3 8500 44900 8700 45000 0 FreeSans 400 0 0 0 a[2]
port 5 nsew signal input
flabel metal3 9100 44900 9300 45000 0 FreeSans 400 0 0 0 a[3]
port 6 nsew signal input
flabel metal3 9700 44900 9900 45000 0 FreeSans 400 0 0 0 a[4]
port 7 nsew signal input
flabel metal3 10300 44900 10500 45000 0 FreeSans 400 0 0 0 a[5]
port 8 nsew signal input
flabel metal3 10900 44900 11100 45000 0 FreeSans 400 0 0 0 a[6]
port 9 nsew signal input
flabel metal3 11500 44900 11700 45000 0 FreeSans 400 0 0 0 a[7]
port 10 nsew signal input
flabel metal3 12100 44900 12300 45000 0 FreeSans 400 0 0 0 a[8]
port 11 nsew signal input
flabel metal2 8770 42772 11190 42872 0 FreeSans 320 0 0 0 a[8]
flabel metal2 8770 42634 11190 42734 0 FreeSans 320 0 0 0 a[7]
flabel metal2 8770 42496 11190 42596 0 FreeSans 320 0 0 0 a[6]
flabel metal2 8770 42358 11190 42458 0 FreeSans 320 0 0 0 a[5]
flabel metal2 8770 42220 11190 42320 0 FreeSans 320 0 0 0 a[4]
flabel metal3 8774 42880 8974 42960 0 FreeSans 320 0 0 0 a[0]
flabel metal3 9042 42880 9242 42960 0 FreeSans 320 0 0 0 a[1]
flabel metal3 9310 42880 9510 42960 0 FreeSans 320 0 0 0 a[2]
flabel metal3 9578 42880 9778 42960 0 FreeSans 320 0 0 0 a[3]
flabel metal3 10114 42880 10314 42960 0 FreeSans 320 0 0 0 a[5]
flabel metal3 10382 42880 10582 42960 0 FreeSans 320 0 0 0 a[6]
flabel metal3 10650 42880 10850 42960 0 FreeSans 320 0 0 0 a[7]
flabel metal3 10918 42880 11118 42960 0 FreeSans 320 0 0 0 a[8]
flabel metal3 9846 42880 10046 42960 0 FreeSans 320 0 0 0 a[4]
flabel metal2 3747 41595 3797 41645 0 FreeSans 80 0 0 0 l_row_en[0]
flabel metal2 3747 41195 3797 41245 0 FreeSans 80 0 0 0 l_row_en[1]
flabel metal2 3747 40795 3797 40845 0 FreeSans 80 0 0 0 l_row_en[2]
flabel metal2 3747 40395 3797 40445 0 FreeSans 80 0 0 0 l_row_en[3]
flabel metal2 3747 39995 3797 40045 0 FreeSans 80 0 0 0 l_row_en[4]
flabel metal2 3747 39595 3797 39645 0 FreeSans 80 0 0 0 l_row_en[5]
flabel metal2 3747 39195 3797 39245 0 FreeSans 80 0 0 0 l_row_en[6]
flabel metal2 3747 38795 3797 38845 0 FreeSans 80 0 0 0 l_row_en[7]
flabel metal2 3747 38395 3797 38445 0 FreeSans 80 0 0 0 l_row_en[8]
flabel metal2 3747 37995 3797 38045 0 FreeSans 80 0 0 0 l_row_en[9]
flabel metal2 3747 37595 3797 37645 0 FreeSans 80 0 0 0 l_row_en[10]
flabel metal2 3747 37195 3797 37245 0 FreeSans 80 0 0 0 l_row_en[11]
flabel metal2 3747 36795 3797 36845 0 FreeSans 80 0 0 0 l_row_en[12]
flabel metal2 3747 36395 3797 36445 0 FreeSans 80 0 0 0 l_row_en[13]
flabel metal2 3747 35995 3797 36045 0 FreeSans 80 0 0 0 l_row_en[14]
flabel metal2 3747 35595 3797 35645 0 FreeSans 80 0 0 0 l_row_en[15]
flabel metal2 3747 35195 3797 35245 0 FreeSans 80 0 0 0 l_row_en[16]
flabel metal2 3747 34795 3797 34845 0 FreeSans 80 0 0 0 l_row_en[17]
flabel metal2 3747 34395 3797 34445 0 FreeSans 80 0 0 0 l_row_en[18]
flabel metal2 3747 33995 3797 34045 0 FreeSans 80 0 0 0 l_row_en[19]
flabel metal2 3747 33595 3797 33645 0 FreeSans 80 0 0 0 l_row_en[20]
flabel metal2 3747 33195 3797 33245 0 FreeSans 80 0 0 0 l_row_en[21]
flabel metal2 3747 32795 3797 32845 0 FreeSans 80 0 0 0 l_row_en[22]
flabel metal2 3747 32395 3797 32445 0 FreeSans 80 0 0 0 l_row_en[23]
flabel metal2 3747 31995 3797 32045 0 FreeSans 80 0 0 0 l_row_en[24]
flabel metal2 3747 31595 3797 31645 0 FreeSans 80 0 0 0 l_row_en[25]
flabel metal2 3747 31195 3797 31245 0 FreeSans 80 0 0 0 l_row_en[26]
flabel metal2 3747 30795 3797 30845 0 FreeSans 80 0 0 0 l_row_en[27]
flabel metal2 3747 30395 3797 30445 0 FreeSans 80 0 0 0 l_row_en[28]
flabel metal2 3747 29995 3797 30045 0 FreeSans 80 0 0 0 l_row_en[29]
flabel metal2 3747 29595 3797 29645 0 FreeSans 80 0 0 0 l_row_en[30]
flabel metal2 3747 29195 3797 29245 0 FreeSans 80 0 0 0 l_row_en[31]
flabel metal2 3747 41531 3797 41581 0 FreeSans 80 0 0 0 l_row_en_b[0]
flabel metal2 3747 41131 3797 41181 0 FreeSans 80 0 0 0 l_row_en_b[1]
flabel metal2 3747 40731 3797 40781 0 FreeSans 80 0 0 0 l_row_en_b[2]
flabel metal2 3747 40331 3797 40381 0 FreeSans 80 0 0 0 l_row_en_b[3]
flabel metal2 3747 39931 3797 39981 0 FreeSans 80 0 0 0 l_row_en_b[4]
flabel metal2 3747 39531 3797 39581 0 FreeSans 80 0 0 0 l_row_en_b[5]
flabel metal2 3747 39131 3797 39181 0 FreeSans 80 0 0 0 l_row_en_b[6]
flabel metal2 3747 38731 3797 38781 0 FreeSans 80 0 0 0 l_row_en_b[7]
flabel metal2 3747 38331 3797 38381 0 FreeSans 80 0 0 0 l_row_en_b[8]
flabel metal2 3747 37931 3797 37981 0 FreeSans 80 0 0 0 l_row_en_b[9]
flabel metal2 3747 37531 3797 37581 0 FreeSans 80 0 0 0 l_row_en_b[10]
flabel metal2 3747 37131 3797 37181 0 FreeSans 80 0 0 0 l_row_en_b[11]
flabel metal2 3747 36731 3797 36781 0 FreeSans 80 0 0 0 l_row_en_b[12]
flabel metal2 3747 36331 3797 36381 0 FreeSans 80 0 0 0 l_row_en_b[13]
flabel metal2 3747 35931 3797 35981 0 FreeSans 80 0 0 0 l_row_en_b[14]
flabel metal2 3747 35531 3797 35581 0 FreeSans 80 0 0 0 l_row_en_b[15]
flabel metal2 3747 35131 3797 35181 0 FreeSans 80 0 0 0 l_row_en_b[16]
flabel metal2 3747 34731 3797 34781 0 FreeSans 80 0 0 0 l_row_en_b[17]
flabel metal2 3747 34331 3797 34381 0 FreeSans 80 0 0 0 l_row_en_b[18]
flabel metal2 3747 33931 3797 33981 0 FreeSans 80 0 0 0 l_row_en_b[19]
flabel metal2 3747 33531 3797 33581 0 FreeSans 80 0 0 0 l_row_en_b[20]
flabel metal2 3747 33131 3797 33181 0 FreeSans 80 0 0 0 l_row_en_b[21]
flabel metal2 3747 32731 3797 32781 0 FreeSans 80 0 0 0 l_row_en_b[22]
flabel metal2 3747 32331 3797 32381 0 FreeSans 80 0 0 0 l_row_en_b[23]
flabel metal2 3747 31931 3797 31981 0 FreeSans 80 0 0 0 l_row_en_b[24]
flabel metal2 3747 31531 3797 31581 0 FreeSans 80 0 0 0 l_row_en_b[25]
flabel metal2 3747 31131 3797 31181 0 FreeSans 80 0 0 0 l_row_en_b[26]
flabel metal2 3747 30731 3797 30781 0 FreeSans 80 0 0 0 l_row_en_b[27]
flabel metal2 3747 30331 3797 30381 0 FreeSans 80 0 0 0 l_row_en_b[28]
flabel metal2 3747 29931 3797 29981 0 FreeSans 80 0 0 0 l_row_en_b[29]
flabel metal2 3747 29531 3797 29581 0 FreeSans 80 0 0 0 l_row_en_b[30]
flabel metal2 3747 29131 3797 29181 0 FreeSans 80 0 0 0 l_row_en_b[31]
flabel metal2 16163 41595 16213 41645 0 FreeSans 80 0 0 0 r_row_en[0]
flabel metal2 16163 41195 16213 41245 0 FreeSans 80 0 0 0 r_row_en[1]
flabel metal2 16163 40795 16213 40845 0 FreeSans 80 0 0 0 r_row_en[2]
flabel metal2 16163 40395 16213 40445 0 FreeSans 80 0 0 0 r_row_en[3]
flabel metal2 16163 39995 16213 40045 0 FreeSans 80 0 0 0 r_row_en[4]
flabel metal2 16163 39595 16213 39645 0 FreeSans 80 0 0 0 r_row_en[5]
flabel metal2 16163 39195 16213 39245 0 FreeSans 80 0 0 0 r_row_en[6]
flabel metal2 16163 38795 16213 38845 0 FreeSans 80 0 0 0 r_row_en[7]
flabel metal2 16163 38395 16213 38445 0 FreeSans 80 0 0 0 r_row_en[8]
flabel metal2 16163 37995 16213 38045 0 FreeSans 80 0 0 0 r_row_en[9]
flabel metal2 16163 37595 16213 37645 0 FreeSans 80 0 0 0 r_row_en[10]
flabel metal2 16163 37195 16213 37245 0 FreeSans 80 0 0 0 r_row_en[11]
flabel metal2 16163 36795 16213 36845 0 FreeSans 80 0 0 0 r_row_en[12]
flabel metal2 16163 36395 16213 36445 0 FreeSans 80 0 0 0 r_row_en[13]
flabel metal2 16163 35995 16213 36045 0 FreeSans 80 0 0 0 r_row_en[14]
flabel metal2 16163 35595 16213 35645 0 FreeSans 80 0 0 0 r_row_en[15]
flabel metal2 16163 35195 16213 35245 0 FreeSans 80 0 0 0 r_row_en[16]
flabel metal2 16163 34795 16213 34845 0 FreeSans 80 0 0 0 r_row_en[17]
flabel metal2 16163 34395 16213 34445 0 FreeSans 80 0 0 0 r_row_en[18]
flabel metal2 16163 33995 16213 34045 0 FreeSans 80 0 0 0 r_row_en[19]
flabel metal2 16163 33595 16213 33645 0 FreeSans 80 0 0 0 r_row_en[20]
flabel metal2 16163 33195 16213 33245 0 FreeSans 80 0 0 0 r_row_en[21]
flabel metal2 16163 32795 16213 32845 0 FreeSans 80 0 0 0 r_row_en[22]
flabel metal2 16163 32395 16213 32445 0 FreeSans 80 0 0 0 r_row_en[23]
flabel metal2 16163 31995 16213 32045 0 FreeSans 80 0 0 0 r_row_en[24]
flabel metal2 16163 31595 16213 31645 0 FreeSans 80 0 0 0 r_row_en[25]
flabel metal2 16163 31195 16213 31245 0 FreeSans 80 0 0 0 r_row_en[26]
flabel metal2 16163 30795 16213 30845 0 FreeSans 80 0 0 0 r_row_en[27]
flabel metal2 16163 30395 16213 30445 0 FreeSans 80 0 0 0 r_row_en[28]
flabel metal2 16163 29995 16213 30045 0 FreeSans 80 0 0 0 r_row_en[29]
flabel metal2 16163 29595 16213 29645 0 FreeSans 80 0 0 0 r_row_en[30]
flabel metal2 16163 29195 16213 29245 0 FreeSans 80 0 0 0 r_row_en[31]
flabel metal2 16163 41531 16213 41581 0 FreeSans 80 0 0 0 r_row_en_b[0]
flabel metal2 16163 41131 16213 41181 0 FreeSans 80 0 0 0 r_row_en_b[1]
flabel metal2 16163 40731 16213 40781 0 FreeSans 80 0 0 0 r_row_en_b[2]
flabel metal2 16163 40331 16213 40381 0 FreeSans 80 0 0 0 r_row_en_b[3]
flabel metal2 16163 39931 16213 39981 0 FreeSans 80 0 0 0 r_row_en_b[4]
flabel metal2 16163 39531 16213 39581 0 FreeSans 80 0 0 0 r_row_en_b[5]
flabel metal2 16163 39131 16213 39181 0 FreeSans 80 0 0 0 r_row_en_b[6]
flabel metal2 16163 38731 16213 38781 0 FreeSans 80 0 0 0 r_row_en_b[7]
flabel metal2 16163 38331 16213 38381 0 FreeSans 80 0 0 0 r_row_en_b[8]
flabel metal2 16163 37931 16213 37981 0 FreeSans 80 0 0 0 r_row_en_b[9]
flabel metal2 16163 37531 16213 37581 0 FreeSans 80 0 0 0 r_row_en_b[10]
flabel metal2 16163 37131 16213 37181 0 FreeSans 80 0 0 0 r_row_en_b[11]
flabel metal2 16163 36731 16213 36781 0 FreeSans 80 0 0 0 r_row_en_b[12]
flabel metal2 16163 36331 16213 36381 0 FreeSans 80 0 0 0 r_row_en_b[13]
flabel metal2 16163 35931 16213 35981 0 FreeSans 80 0 0 0 r_row_en_b[14]
flabel metal2 16163 35531 16213 35581 0 FreeSans 80 0 0 0 r_row_en_b[15]
flabel metal2 16163 35131 16213 35181 0 FreeSans 80 0 0 0 r_row_en_b[16]
flabel metal2 16163 34731 16213 34781 0 FreeSans 80 0 0 0 r_row_en_b[17]
flabel metal2 16163 34331 16213 34381 0 FreeSans 80 0 0 0 r_row_en_b[18]
flabel metal2 16163 33931 16213 33981 0 FreeSans 80 0 0 0 r_row_en_b[19]
flabel metal2 16163 33531 16213 33581 0 FreeSans 80 0 0 0 r_row_en_b[20]
flabel metal2 16163 33131 16213 33181 0 FreeSans 80 0 0 0 r_row_en_b[21]
flabel metal2 16163 32731 16213 32781 0 FreeSans 80 0 0 0 r_row_en_b[22]
flabel metal2 16163 32331 16213 32381 0 FreeSans 80 0 0 0 r_row_en_b[23]
flabel metal2 16163 31931 16213 31981 0 FreeSans 80 0 0 0 r_row_en_b[24]
flabel metal2 16163 31531 16213 31581 0 FreeSans 80 0 0 0 r_row_en_b[25]
flabel metal2 16163 31131 16213 31181 0 FreeSans 80 0 0 0 r_row_en_b[26]
flabel metal2 16163 30731 16213 30781 0 FreeSans 80 0 0 0 r_row_en_b[27]
flabel metal2 16163 30331 16213 30381 0 FreeSans 80 0 0 0 r_row_en_b[28]
flabel metal2 16163 29931 16213 29981 0 FreeSans 80 0 0 0 r_row_en_b[29]
flabel metal2 16163 29531 16213 29581 0 FreeSans 80 0 0 0 r_row_en_b[30]
flabel metal2 16163 29131 16213 29181 0 FreeSans 80 0 0 0 r_row_en_b[31]
flabel metal3 5100 44900 5900 45000 0 FreeSans 400 0 0 0 VPWR
port 1 nsew power default
flabel metal3 12700 44900 13500 45000 0 FreeSans 400 0 0 0 VPWR
port 1 nsew power default
flabel metal3 6100 44900 6900 45000 0 FreeSans 400 0 0 0 VGND
port 2 nsew ground default
flabel metal3 13700 44900 14500 45000 0 FreeSans 400 0 0 0 VGND
port 2 nsew ground default
flabel metal2 4989 41532 5047 41590 0 FreeSans 160 0 0 0 l_w[0]
flabel metal2 4989 41132 5047 41190 0 FreeSans 160 0 0 0 l_w[1]
flabel metal2 4989 40732 5047 40790 0 FreeSans 160 0 0 0 l_w[2]
flabel metal2 4989 40332 5047 40390 0 FreeSans 160 0 0 0 l_w[3]
flabel metal2 4989 39932 5047 39990 0 FreeSans 160 0 0 0 l_w[4]
flabel metal2 4989 39532 5047 39590 0 FreeSans 160 0 0 0 l_w[5]
flabel metal2 4989 39132 5047 39190 0 FreeSans 160 0 0 0 l_w[6]
flabel metal2 4989 38732 5047 38790 0 FreeSans 160 0 0 0 l_w[7]
flabel metal2 4989 38332 5047 38390 0 FreeSans 160 0 0 0 l_w[8]
flabel metal2 4989 37932 5047 37990 0 FreeSans 160 0 0 0 l_w[9]
flabel metal2 4989 37532 5047 37590 0 FreeSans 160 0 0 0 l_w[10]
flabel metal2 4989 37132 5047 37190 0 FreeSans 160 0 0 0 l_w[11]
flabel metal2 4989 36732 5047 36790 0 FreeSans 160 0 0 0 l_w[12]
flabel metal2 4989 36332 5047 36390 0 FreeSans 160 0 0 0 l_w[13]
flabel metal2 4989 35932 5047 35990 0 FreeSans 160 0 0 0 l_w[14]
flabel metal2 4989 35532 5047 35590 0 FreeSans 160 0 0 0 l_w[15]
flabel metal2 4989 35132 5047 35190 0 FreeSans 160 0 0 0 l_w[16]
flabel metal2 4989 34732 5047 34790 0 FreeSans 160 0 0 0 l_w[17]
flabel metal2 4989 34332 5047 34390 0 FreeSans 160 0 0 0 l_w[18]
flabel metal2 4989 33932 5047 33990 0 FreeSans 160 0 0 0 l_w[19]
flabel metal2 4989 33532 5047 33590 0 FreeSans 160 0 0 0 l_w[20]
flabel metal2 4989 33132 5047 33190 0 FreeSans 160 0 0 0 l_w[21]
flabel metal2 4989 32732 5047 32790 0 FreeSans 160 0 0 0 l_w[22]
flabel metal2 4989 32332 5047 32390 0 FreeSans 160 0 0 0 l_w[23]
flabel metal2 4989 31932 5047 31990 0 FreeSans 160 0 0 0 l_w[24]
flabel metal2 4989 31532 5047 31590 0 FreeSans 160 0 0 0 l_w[25]
flabel metal2 4989 31132 5047 31190 0 FreeSans 160 0 0 0 l_w[26]
flabel metal2 4989 30732 5047 30790 0 FreeSans 160 0 0 0 l_w[27]
flabel metal2 4989 30332 5047 30390 0 FreeSans 160 0 0 0 l_w[28]
flabel metal2 4989 29932 5047 29990 0 FreeSans 160 0 0 0 l_w[29]
flabel metal2 4989 29532 5047 29590 0 FreeSans 160 0 0 0 l_w[30]
flabel metal2 4989 29132 5047 29190 0 FreeSans 160 0 0 0 l_w[31]
flabel metal2 14913 41532 14971 41590 0 FreeSans 160 0 0 0 r_w[0]
flabel metal2 14913 41132 14971 41190 0 FreeSans 160 0 0 0 r_w[1]
flabel metal2 14913 40732 14971 40790 0 FreeSans 160 0 0 0 r_w[2]
flabel metal2 14913 40332 14971 40390 0 FreeSans 160 0 0 0 r_w[3]
flabel metal2 14913 39932 14971 39990 0 FreeSans 160 0 0 0 r_w[4]
flabel metal2 14913 39532 14971 39590 0 FreeSans 160 0 0 0 r_w[5]
flabel metal2 14913 39132 14971 39190 0 FreeSans 160 0 0 0 r_w[6]
flabel metal2 14913 38732 14971 38790 0 FreeSans 160 0 0 0 r_w[7]
flabel metal2 14913 38332 14971 38390 0 FreeSans 160 0 0 0 r_w[8]
flabel metal2 14913 37932 14971 37990 0 FreeSans 160 0 0 0 r_w[9]
flabel metal2 14913 37532 14971 37590 0 FreeSans 160 0 0 0 r_w[10]
flabel metal2 14913 37132 14971 37190 0 FreeSans 160 0 0 0 r_w[11]
flabel metal2 14913 36732 14971 36790 0 FreeSans 160 0 0 0 r_w[12]
flabel metal2 14913 36332 14971 36390 0 FreeSans 160 0 0 0 r_w[13]
flabel metal2 14913 35932 14971 35990 0 FreeSans 160 0 0 0 r_w[14]
flabel metal2 14913 35532 14971 35590 0 FreeSans 160 0 0 0 r_w[15]
flabel metal2 14913 35132 14971 35190 0 FreeSans 160 0 0 0 r_w[16]
flabel metal2 14913 34732 14971 34790 0 FreeSans 160 0 0 0 r_w[17]
flabel metal2 14913 34332 14971 34390 0 FreeSans 160 0 0 0 r_w[18]
flabel metal2 14913 33932 14971 33990 0 FreeSans 160 0 0 0 r_w[19]
flabel metal2 14913 33532 14971 33590 0 FreeSans 160 0 0 0 r_w[20]
flabel metal2 14913 33132 14971 33190 0 FreeSans 160 0 0 0 r_w[21]
flabel metal2 14913 32732 14971 32790 0 FreeSans 160 0 0 0 r_w[22]
flabel metal2 14913 32332 14971 32390 0 FreeSans 160 0 0 0 r_w[23]
flabel metal2 14913 31932 14971 31990 0 FreeSans 160 0 0 0 r_w[24]
flabel metal2 14913 31532 14971 31590 0 FreeSans 160 0 0 0 r_w[25]
flabel metal2 14913 31132 14971 31190 0 FreeSans 160 0 0 0 r_w[26]
flabel metal2 14913 30732 14971 30790 0 FreeSans 160 0 0 0 r_w[27]
flabel metal2 14913 30332 14971 30390 0 FreeSans 160 0 0 0 r_w[28]
flabel metal2 14913 29932 14971 29990 0 FreeSans 160 0 0 0 r_w[29]
flabel metal2 14913 29532 14971 29590 0 FreeSans 160 0 0 0 r_w[30]
flabel metal2 14913 29132 14971 29190 0 FreeSans 160 0 0 0 r_w[31]
flabel metal5 -19900 -1400 38500 -600 0 FreeSans 3200 0 0 0 VTUN
<< end >>
