magic
tech sky130A
timestamp 1716993426
<< checkpaint >>
rect -652 -630 994 870
use fgcell_amp  x1
timestamp 1716993254
transform 1 0 0 0 1 3000
box 0 -3000 101 100
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC1
timestamp 0
transform 1 0 171 0 1 120
box -193 -120 193 120
<< end >>
