magic
tech sky130A
timestamp 1717164252
<< error_p >>
rect 349 5374 580 5454
rect 2349 5374 2580 5454
rect 4349 5374 4580 5454
rect 6349 5374 6580 5454
rect 8349 5374 8580 5454
rect 10349 5374 10580 5454
rect 12349 5374 12580 5454
rect 14349 5374 14580 5454
rect 16349 5374 16580 5454
rect 18349 5374 18580 5454
rect 349 3874 580 3954
rect 2349 3874 2580 3954
rect 4349 3874 4580 3954
rect 6349 3874 6580 3954
rect 8349 3874 8580 3954
rect 10349 3874 10580 3954
rect 12349 3874 12580 3954
rect 14349 3874 14580 3954
rect 16349 3874 16580 3954
rect 18349 3874 18580 3954
rect 349 2374 580 2454
rect 2349 2374 2580 2454
rect 4349 2374 4580 2454
rect 6349 2374 6580 2454
rect 8349 2374 8580 2454
rect 10349 2374 10580 2454
rect 12349 2374 12580 2454
rect 14349 2374 14580 2454
rect 16349 2374 16580 2454
rect 18349 2374 18580 2454
rect 349 874 580 954
rect 2349 874 2580 954
rect 4349 874 4580 954
rect 6349 874 6580 954
rect 8349 874 8580 954
rect 10349 874 10580 954
rect 12349 874 12580 954
rect 14349 874 14580 954
rect 16349 874 16580 954
rect 18349 874 18580 954
use fgcell_amp_MOS_cap_thick_poly  fgcell_amp_MOS_cap_thick_poly_0
array 0 9 2000 0 4 1500
timestamp 1717163667
transform 1 0 -70 0 1 11105
box 70 -3605 2053 -2482
use fgcell_amp_MOS_cap_thin_poly  fgcell_amp_MOS_cap_thin_poly_0
array 0 9 2000 0 4 1500
timestamp 1717163634
transform 1 0 -70 0 1 3605
box 37 -3605 2053 -2482
<< end >>
