magic
tech sky130A
magscale 1 2
timestamp 1717597427
<< error_p >>
rect 2240 29596 2480 29620
rect 2240 29536 2264 29596
rect 2456 29536 2480 29596
rect 2240 29380 2480 29536
rect 6240 29596 6480 29620
rect 6240 29536 6264 29596
rect 6456 29536 6480 29596
rect 6240 29380 6480 29536
rect 10240 29596 10480 29620
rect 10240 29536 10264 29596
rect 10456 29536 10480 29596
rect 10240 29380 10480 29536
rect 14240 29596 14480 29620
rect 14240 29536 14264 29596
rect 14456 29536 14480 29596
rect 14240 29380 14480 29536
rect 18240 29596 18480 29620
rect 18240 29536 18264 29596
rect 18456 29536 18480 29596
rect 18240 29380 18480 29536
rect 22240 29596 22480 29620
rect 22240 29536 22264 29596
rect 22456 29536 22480 29596
rect 22240 29380 22480 29536
rect 26240 29596 26480 29620
rect 26240 29536 26264 29596
rect 26456 29536 26480 29596
rect 26240 29380 26480 29536
rect 30240 29596 30480 29620
rect 30240 29536 30264 29596
rect 30456 29536 30480 29596
rect 30240 29380 30480 29536
rect 34240 29596 34480 29620
rect 34240 29536 34264 29596
rect 34456 29536 34480 29596
rect 34240 29380 34480 29536
rect 38240 29596 38480 29620
rect 38240 29536 38264 29596
rect 38456 29536 38480 29596
rect 38240 29380 38480 29536
rect 1936 29160 2256 29216
rect 360 28916 600 28940
rect 360 28724 384 28916
rect 576 28724 600 28916
rect 1936 28920 1960 29160
rect 2224 28920 2256 29160
rect 3602 29163 3690 29168
rect 3602 29085 3607 29163
rect 3685 29085 3690 29163
rect 3602 29080 3690 29085
rect 5936 29160 6256 29216
rect 1936 28896 2256 28920
rect 4360 28916 4600 28940
rect 360 28700 600 28724
rect 4360 28724 4384 28916
rect 4576 28724 4600 28916
rect 5936 28920 5960 29160
rect 6224 28920 6256 29160
rect 7602 29163 7690 29168
rect 7602 29085 7607 29163
rect 7685 29085 7690 29163
rect 7602 29080 7690 29085
rect 9936 29160 10256 29216
rect 5936 28896 6256 28920
rect 8360 28916 8600 28940
rect 2810 28711 2946 28716
rect 2810 28637 2815 28711
rect 2941 28637 2946 28711
rect 4360 28700 4600 28724
rect 8360 28724 8384 28916
rect 8576 28724 8600 28916
rect 9936 28920 9960 29160
rect 10224 28920 10256 29160
rect 11602 29163 11690 29168
rect 11602 29085 11607 29163
rect 11685 29085 11690 29163
rect 11602 29080 11690 29085
rect 13936 29160 14256 29216
rect 9936 28896 10256 28920
rect 12360 28916 12600 28940
rect 6810 28711 6946 28716
rect 2810 28632 2946 28637
rect 6810 28637 6815 28711
rect 6941 28637 6946 28711
rect 8360 28700 8600 28724
rect 12360 28724 12384 28916
rect 12576 28724 12600 28916
rect 13936 28920 13960 29160
rect 14224 28920 14256 29160
rect 15602 29163 15690 29168
rect 15602 29085 15607 29163
rect 15685 29085 15690 29163
rect 15602 29080 15690 29085
rect 17936 29160 18256 29216
rect 13936 28896 14256 28920
rect 16360 28916 16600 28940
rect 10810 28711 10946 28716
rect 6810 28632 6946 28637
rect 10810 28637 10815 28711
rect 10941 28637 10946 28711
rect 12360 28700 12600 28724
rect 16360 28724 16384 28916
rect 16576 28724 16600 28916
rect 17936 28920 17960 29160
rect 18224 28920 18256 29160
rect 19602 29163 19690 29168
rect 19602 29085 19607 29163
rect 19685 29085 19690 29163
rect 19602 29080 19690 29085
rect 21936 29160 22256 29216
rect 17936 28896 18256 28920
rect 20360 28916 20600 28940
rect 14810 28711 14946 28716
rect 10810 28632 10946 28637
rect 14810 28637 14815 28711
rect 14941 28637 14946 28711
rect 16360 28700 16600 28724
rect 20360 28724 20384 28916
rect 20576 28724 20600 28916
rect 21936 28920 21960 29160
rect 22224 28920 22256 29160
rect 23602 29163 23690 29168
rect 23602 29085 23607 29163
rect 23685 29085 23690 29163
rect 23602 29080 23690 29085
rect 25936 29160 26256 29216
rect 21936 28896 22256 28920
rect 24360 28916 24600 28940
rect 18810 28711 18946 28716
rect 14810 28632 14946 28637
rect 18810 28637 18815 28711
rect 18941 28637 18946 28711
rect 20360 28700 20600 28724
rect 24360 28724 24384 28916
rect 24576 28724 24600 28916
rect 25936 28920 25960 29160
rect 26224 28920 26256 29160
rect 27602 29163 27690 29168
rect 27602 29085 27607 29163
rect 27685 29085 27690 29163
rect 27602 29080 27690 29085
rect 29936 29160 30256 29216
rect 25936 28896 26256 28920
rect 28360 28916 28600 28940
rect 22810 28711 22946 28716
rect 18810 28632 18946 28637
rect 22810 28637 22815 28711
rect 22941 28637 22946 28711
rect 24360 28700 24600 28724
rect 28360 28724 28384 28916
rect 28576 28724 28600 28916
rect 29936 28920 29960 29160
rect 30224 28920 30256 29160
rect 31602 29163 31690 29168
rect 31602 29085 31607 29163
rect 31685 29085 31690 29163
rect 31602 29080 31690 29085
rect 33936 29160 34256 29216
rect 29936 28896 30256 28920
rect 32360 28916 32600 28940
rect 26810 28711 26946 28716
rect 22810 28632 22946 28637
rect 26810 28637 26815 28711
rect 26941 28637 26946 28711
rect 28360 28700 28600 28724
rect 32360 28724 32384 28916
rect 32576 28724 32600 28916
rect 33936 28920 33960 29160
rect 34224 28920 34256 29160
rect 35602 29163 35690 29168
rect 35602 29085 35607 29163
rect 35685 29085 35690 29163
rect 35602 29080 35690 29085
rect 37936 29160 38256 29216
rect 33936 28896 34256 28920
rect 36360 28916 36600 28940
rect 30810 28711 30946 28716
rect 26810 28632 26946 28637
rect 30810 28637 30815 28711
rect 30941 28637 30946 28711
rect 32360 28700 32600 28724
rect 36360 28724 36384 28916
rect 36576 28724 36600 28916
rect 37936 28920 37960 29160
rect 38224 28920 38256 29160
rect 39602 29163 39690 29168
rect 39602 29085 39607 29163
rect 39685 29085 39690 29163
rect 39602 29080 39690 29085
rect 37936 28896 38256 28920
rect 34810 28711 34946 28716
rect 30810 28632 30946 28637
rect 34810 28637 34815 28711
rect 34941 28637 34946 28711
rect 36360 28700 36600 28724
rect 38810 28711 38946 28716
rect 34810 28632 34946 28637
rect 38810 28637 38815 28711
rect 38941 28637 38946 28711
rect 38810 28632 38946 28637
rect 2338 28573 2518 28574
rect 2338 28395 2339 28573
rect 2517 28395 2518 28573
rect 2338 28394 2518 28395
rect 6338 28573 6518 28574
rect 6338 28395 6339 28573
rect 6517 28395 6518 28573
rect 6338 28394 6518 28395
rect 10338 28573 10518 28574
rect 10338 28395 10339 28573
rect 10517 28395 10518 28573
rect 10338 28394 10518 28395
rect 14338 28573 14518 28574
rect 14338 28395 14339 28573
rect 14517 28395 14518 28573
rect 14338 28394 14518 28395
rect 18338 28573 18518 28574
rect 18338 28395 18339 28573
rect 18517 28395 18518 28573
rect 18338 28394 18518 28395
rect 22338 28573 22518 28574
rect 22338 28395 22339 28573
rect 22517 28395 22518 28573
rect 22338 28394 22518 28395
rect 26338 28573 26518 28574
rect 26338 28395 26339 28573
rect 26517 28395 26518 28573
rect 26338 28394 26518 28395
rect 30338 28573 30518 28574
rect 30338 28395 30339 28573
rect 30517 28395 30518 28573
rect 30338 28394 30518 28395
rect 34338 28573 34518 28574
rect 34338 28395 34339 28573
rect 34517 28395 34518 28573
rect 34338 28394 34518 28395
rect 38338 28573 38518 28574
rect 38338 28395 38339 28573
rect 38517 28395 38518 28573
rect 38338 28394 38518 28395
rect 400 27999 580 28000
rect 400 27821 401 27999
rect 579 27821 580 27999
rect 3734 27996 3740 28002
rect 3780 27996 3786 28002
rect 4400 27999 4580 28000
rect 3728 27990 3734 27996
rect 3786 27990 3792 27996
rect 3728 27944 3734 27950
rect 3786 27944 3792 27950
rect 3734 27938 3740 27944
rect 3780 27938 3786 27944
rect 400 27820 580 27821
rect 4400 27821 4401 27999
rect 4579 27821 4580 27999
rect 7734 27996 7740 28002
rect 7780 27996 7786 28002
rect 8400 27999 8580 28000
rect 7728 27990 7734 27996
rect 7786 27990 7792 27996
rect 7728 27944 7734 27950
rect 7786 27944 7792 27950
rect 7734 27938 7740 27944
rect 7780 27938 7786 27944
rect 4400 27820 4580 27821
rect 8400 27821 8401 27999
rect 8579 27821 8580 27999
rect 11734 27996 11740 28002
rect 11780 27996 11786 28002
rect 12400 27999 12580 28000
rect 11728 27990 11734 27996
rect 11786 27990 11792 27996
rect 11728 27944 11734 27950
rect 11786 27944 11792 27950
rect 11734 27938 11740 27944
rect 11780 27938 11786 27944
rect 8400 27820 8580 27821
rect 12400 27821 12401 27999
rect 12579 27821 12580 27999
rect 15734 27996 15740 28002
rect 15780 27996 15786 28002
rect 16400 27999 16580 28000
rect 15728 27990 15734 27996
rect 15786 27990 15792 27996
rect 15728 27944 15734 27950
rect 15786 27944 15792 27950
rect 15734 27938 15740 27944
rect 15780 27938 15786 27944
rect 12400 27820 12580 27821
rect 16400 27821 16401 27999
rect 16579 27821 16580 27999
rect 19734 27996 19740 28002
rect 19780 27996 19786 28002
rect 20400 27999 20580 28000
rect 19728 27990 19734 27996
rect 19786 27990 19792 27996
rect 19728 27944 19734 27950
rect 19786 27944 19792 27950
rect 19734 27938 19740 27944
rect 19780 27938 19786 27944
rect 16400 27820 16580 27821
rect 20400 27821 20401 27999
rect 20579 27821 20580 27999
rect 23734 27996 23740 28002
rect 23780 27996 23786 28002
rect 24400 27999 24580 28000
rect 23728 27990 23734 27996
rect 23786 27990 23792 27996
rect 23728 27944 23734 27950
rect 23786 27944 23792 27950
rect 23734 27938 23740 27944
rect 23780 27938 23786 27944
rect 20400 27820 20580 27821
rect 24400 27821 24401 27999
rect 24579 27821 24580 27999
rect 27734 27996 27740 28002
rect 27780 27996 27786 28002
rect 28400 27999 28580 28000
rect 27728 27990 27734 27996
rect 27786 27990 27792 27996
rect 27728 27944 27734 27950
rect 27786 27944 27792 27950
rect 27734 27938 27740 27944
rect 27780 27938 27786 27944
rect 24400 27820 24580 27821
rect 28400 27821 28401 27999
rect 28579 27821 28580 27999
rect 31734 27996 31740 28002
rect 31780 27996 31786 28002
rect 32400 27999 32580 28000
rect 31728 27990 31734 27996
rect 31786 27990 31792 27996
rect 31728 27944 31734 27950
rect 31786 27944 31792 27950
rect 31734 27938 31740 27944
rect 31780 27938 31786 27944
rect 28400 27820 28580 27821
rect 32400 27821 32401 27999
rect 32579 27821 32580 27999
rect 35734 27996 35740 28002
rect 35780 27996 35786 28002
rect 36400 27999 36580 28000
rect 35728 27990 35734 27996
rect 35786 27990 35792 27996
rect 35728 27944 35734 27950
rect 35786 27944 35792 27950
rect 35734 27938 35740 27944
rect 35780 27938 35786 27944
rect 32400 27820 32580 27821
rect 36400 27821 36401 27999
rect 36579 27821 36580 27999
rect 39734 27996 39740 28002
rect 39780 27996 39786 28002
rect 39728 27990 39734 27996
rect 39786 27990 39792 27996
rect 39728 27944 39734 27950
rect 39786 27944 39792 27950
rect 39734 27938 39740 27944
rect 39780 27938 39786 27944
rect 36400 27820 36580 27821
rect 3262 27808 3268 27814
rect 3308 27808 3314 27814
rect 7262 27808 7268 27814
rect 7308 27808 7314 27814
rect 11262 27808 11268 27814
rect 11308 27808 11314 27814
rect 15262 27808 15268 27814
rect 15308 27808 15314 27814
rect 19262 27808 19268 27814
rect 19308 27808 19314 27814
rect 23262 27808 23268 27814
rect 23308 27808 23314 27814
rect 27262 27808 27268 27814
rect 27308 27808 27314 27814
rect 31262 27808 31268 27814
rect 31308 27808 31314 27814
rect 35262 27808 35268 27814
rect 35308 27808 35314 27814
rect 39262 27808 39268 27814
rect 39308 27808 39314 27814
rect 3256 27802 3262 27808
rect 3314 27802 3320 27808
rect 7256 27802 7262 27808
rect 7314 27802 7320 27808
rect 11256 27802 11262 27808
rect 11314 27802 11320 27808
rect 15256 27802 15262 27808
rect 15314 27802 15320 27808
rect 19256 27802 19262 27808
rect 19314 27802 19320 27808
rect 23256 27802 23262 27808
rect 23314 27802 23320 27808
rect 27256 27802 27262 27808
rect 27314 27802 27320 27808
rect 31256 27802 31262 27808
rect 31314 27802 31320 27808
rect 35256 27802 35262 27808
rect 35314 27802 35320 27808
rect 39256 27802 39262 27808
rect 39314 27802 39320 27808
rect 3256 27756 3262 27762
rect 3314 27756 3320 27762
rect 7256 27756 7262 27762
rect 7314 27756 7320 27762
rect 11256 27756 11262 27762
rect 11314 27756 11320 27762
rect 15256 27756 15262 27762
rect 15314 27756 15320 27762
rect 19256 27756 19262 27762
rect 19314 27756 19320 27762
rect 23256 27756 23262 27762
rect 23314 27756 23320 27762
rect 27256 27756 27262 27762
rect 27314 27756 27320 27762
rect 31256 27756 31262 27762
rect 31314 27756 31320 27762
rect 35256 27756 35262 27762
rect 35314 27756 35320 27762
rect 39256 27756 39262 27762
rect 39314 27756 39320 27762
rect 3262 27750 3268 27756
rect 3308 27750 3314 27756
rect 7262 27750 7268 27756
rect 7308 27750 7314 27756
rect 11262 27750 11268 27756
rect 11308 27750 11314 27756
rect 15262 27750 15268 27756
rect 15308 27750 15314 27756
rect 19262 27750 19268 27756
rect 19308 27750 19314 27756
rect 23262 27750 23268 27756
rect 23308 27750 23314 27756
rect 27262 27750 27268 27756
rect 27308 27750 27314 27756
rect 31262 27750 31268 27756
rect 31308 27750 31314 27756
rect 35262 27750 35268 27756
rect 35308 27750 35314 27756
rect 39262 27750 39268 27756
rect 39308 27750 39314 27756
rect 2240 27296 2480 27320
rect 2240 27104 2264 27296
rect 2456 27104 2480 27296
rect 2240 27080 2480 27104
rect 6240 27296 6480 27320
rect 6240 27104 6264 27296
rect 6456 27104 6480 27296
rect 6240 27080 6480 27104
rect 10240 27296 10480 27320
rect 10240 27104 10264 27296
rect 10456 27104 10480 27296
rect 10240 27080 10480 27104
rect 14240 27296 14480 27320
rect 14240 27104 14264 27296
rect 14456 27104 14480 27296
rect 14240 27080 14480 27104
rect 18240 27296 18480 27320
rect 18240 27104 18264 27296
rect 18456 27104 18480 27296
rect 18240 27080 18480 27104
rect 22240 27296 22480 27320
rect 22240 27104 22264 27296
rect 22456 27104 22480 27296
rect 22240 27080 22480 27104
rect 26240 27296 26480 27320
rect 26240 27104 26264 27296
rect 26456 27104 26480 27296
rect 26240 27080 26480 27104
rect 30240 27296 30480 27320
rect 30240 27104 30264 27296
rect 30456 27104 30480 27296
rect 30240 27080 30480 27104
rect 34240 27296 34480 27320
rect 34240 27104 34264 27296
rect 34456 27104 34480 27296
rect 34240 27080 34480 27104
rect 38240 27296 38480 27320
rect 38240 27104 38264 27296
rect 38456 27104 38480 27296
rect 38240 27080 38480 27104
rect 2240 26596 2480 26620
rect 2240 26536 2264 26596
rect 2456 26536 2480 26596
rect 2240 26380 2480 26536
rect 6240 26596 6480 26620
rect 6240 26536 6264 26596
rect 6456 26536 6480 26596
rect 6240 26380 6480 26536
rect 10240 26596 10480 26620
rect 10240 26536 10264 26596
rect 10456 26536 10480 26596
rect 10240 26380 10480 26536
rect 14240 26596 14480 26620
rect 14240 26536 14264 26596
rect 14456 26536 14480 26596
rect 14240 26380 14480 26536
rect 18240 26596 18480 26620
rect 18240 26536 18264 26596
rect 18456 26536 18480 26596
rect 18240 26380 18480 26536
rect 22240 26596 22480 26620
rect 22240 26536 22264 26596
rect 22456 26536 22480 26596
rect 22240 26380 22480 26536
rect 26240 26596 26480 26620
rect 26240 26536 26264 26596
rect 26456 26536 26480 26596
rect 26240 26380 26480 26536
rect 30240 26596 30480 26620
rect 30240 26536 30264 26596
rect 30456 26536 30480 26596
rect 30240 26380 30480 26536
rect 34240 26596 34480 26620
rect 34240 26536 34264 26596
rect 34456 26536 34480 26596
rect 34240 26380 34480 26536
rect 38240 26596 38480 26620
rect 38240 26536 38264 26596
rect 38456 26536 38480 26596
rect 38240 26380 38480 26536
rect 1936 26160 2256 26216
rect 360 25916 600 25940
rect 360 25724 384 25916
rect 576 25724 600 25916
rect 1936 25920 1960 26160
rect 2224 25920 2256 26160
rect 3602 26163 3690 26168
rect 3602 26085 3607 26163
rect 3685 26085 3690 26163
rect 3602 26080 3690 26085
rect 5936 26160 6256 26216
rect 1936 25896 2256 25920
rect 4360 25916 4600 25940
rect 360 25700 600 25724
rect 4360 25724 4384 25916
rect 4576 25724 4600 25916
rect 5936 25920 5960 26160
rect 6224 25920 6256 26160
rect 7602 26163 7690 26168
rect 7602 26085 7607 26163
rect 7685 26085 7690 26163
rect 7602 26080 7690 26085
rect 9936 26160 10256 26216
rect 5936 25896 6256 25920
rect 8360 25916 8600 25940
rect 2810 25711 2946 25716
rect 2810 25637 2815 25711
rect 2941 25637 2946 25711
rect 4360 25700 4600 25724
rect 8360 25724 8384 25916
rect 8576 25724 8600 25916
rect 9936 25920 9960 26160
rect 10224 25920 10256 26160
rect 11602 26163 11690 26168
rect 11602 26085 11607 26163
rect 11685 26085 11690 26163
rect 11602 26080 11690 26085
rect 13936 26160 14256 26216
rect 9936 25896 10256 25920
rect 12360 25916 12600 25940
rect 6810 25711 6946 25716
rect 2810 25632 2946 25637
rect 6810 25637 6815 25711
rect 6941 25637 6946 25711
rect 8360 25700 8600 25724
rect 12360 25724 12384 25916
rect 12576 25724 12600 25916
rect 13936 25920 13960 26160
rect 14224 25920 14256 26160
rect 15602 26163 15690 26168
rect 15602 26085 15607 26163
rect 15685 26085 15690 26163
rect 15602 26080 15690 26085
rect 17936 26160 18256 26216
rect 13936 25896 14256 25920
rect 16360 25916 16600 25940
rect 10810 25711 10946 25716
rect 6810 25632 6946 25637
rect 10810 25637 10815 25711
rect 10941 25637 10946 25711
rect 12360 25700 12600 25724
rect 16360 25724 16384 25916
rect 16576 25724 16600 25916
rect 17936 25920 17960 26160
rect 18224 25920 18256 26160
rect 19602 26163 19690 26168
rect 19602 26085 19607 26163
rect 19685 26085 19690 26163
rect 19602 26080 19690 26085
rect 21936 26160 22256 26216
rect 17936 25896 18256 25920
rect 20360 25916 20600 25940
rect 14810 25711 14946 25716
rect 10810 25632 10946 25637
rect 14810 25637 14815 25711
rect 14941 25637 14946 25711
rect 16360 25700 16600 25724
rect 20360 25724 20384 25916
rect 20576 25724 20600 25916
rect 21936 25920 21960 26160
rect 22224 25920 22256 26160
rect 23602 26163 23690 26168
rect 23602 26085 23607 26163
rect 23685 26085 23690 26163
rect 23602 26080 23690 26085
rect 25936 26160 26256 26216
rect 21936 25896 22256 25920
rect 24360 25916 24600 25940
rect 18810 25711 18946 25716
rect 14810 25632 14946 25637
rect 18810 25637 18815 25711
rect 18941 25637 18946 25711
rect 20360 25700 20600 25724
rect 24360 25724 24384 25916
rect 24576 25724 24600 25916
rect 25936 25920 25960 26160
rect 26224 25920 26256 26160
rect 27602 26163 27690 26168
rect 27602 26085 27607 26163
rect 27685 26085 27690 26163
rect 27602 26080 27690 26085
rect 29936 26160 30256 26216
rect 25936 25896 26256 25920
rect 28360 25916 28600 25940
rect 22810 25711 22946 25716
rect 18810 25632 18946 25637
rect 22810 25637 22815 25711
rect 22941 25637 22946 25711
rect 24360 25700 24600 25724
rect 28360 25724 28384 25916
rect 28576 25724 28600 25916
rect 29936 25920 29960 26160
rect 30224 25920 30256 26160
rect 31602 26163 31690 26168
rect 31602 26085 31607 26163
rect 31685 26085 31690 26163
rect 31602 26080 31690 26085
rect 33936 26160 34256 26216
rect 29936 25896 30256 25920
rect 32360 25916 32600 25940
rect 26810 25711 26946 25716
rect 22810 25632 22946 25637
rect 26810 25637 26815 25711
rect 26941 25637 26946 25711
rect 28360 25700 28600 25724
rect 32360 25724 32384 25916
rect 32576 25724 32600 25916
rect 33936 25920 33960 26160
rect 34224 25920 34256 26160
rect 35602 26163 35690 26168
rect 35602 26085 35607 26163
rect 35685 26085 35690 26163
rect 35602 26080 35690 26085
rect 37936 26160 38256 26216
rect 33936 25896 34256 25920
rect 36360 25916 36600 25940
rect 30810 25711 30946 25716
rect 26810 25632 26946 25637
rect 30810 25637 30815 25711
rect 30941 25637 30946 25711
rect 32360 25700 32600 25724
rect 36360 25724 36384 25916
rect 36576 25724 36600 25916
rect 37936 25920 37960 26160
rect 38224 25920 38256 26160
rect 39602 26163 39690 26168
rect 39602 26085 39607 26163
rect 39685 26085 39690 26163
rect 39602 26080 39690 26085
rect 37936 25896 38256 25920
rect 34810 25711 34946 25716
rect 30810 25632 30946 25637
rect 34810 25637 34815 25711
rect 34941 25637 34946 25711
rect 36360 25700 36600 25724
rect 38810 25711 38946 25716
rect 34810 25632 34946 25637
rect 38810 25637 38815 25711
rect 38941 25637 38946 25711
rect 38810 25632 38946 25637
rect 2338 25573 2518 25574
rect 2338 25395 2339 25573
rect 2517 25395 2518 25573
rect 2338 25394 2518 25395
rect 6338 25573 6518 25574
rect 6338 25395 6339 25573
rect 6517 25395 6518 25573
rect 6338 25394 6518 25395
rect 10338 25573 10518 25574
rect 10338 25395 10339 25573
rect 10517 25395 10518 25573
rect 10338 25394 10518 25395
rect 14338 25573 14518 25574
rect 14338 25395 14339 25573
rect 14517 25395 14518 25573
rect 14338 25394 14518 25395
rect 18338 25573 18518 25574
rect 18338 25395 18339 25573
rect 18517 25395 18518 25573
rect 18338 25394 18518 25395
rect 22338 25573 22518 25574
rect 22338 25395 22339 25573
rect 22517 25395 22518 25573
rect 22338 25394 22518 25395
rect 26338 25573 26518 25574
rect 26338 25395 26339 25573
rect 26517 25395 26518 25573
rect 26338 25394 26518 25395
rect 30338 25573 30518 25574
rect 30338 25395 30339 25573
rect 30517 25395 30518 25573
rect 30338 25394 30518 25395
rect 34338 25573 34518 25574
rect 34338 25395 34339 25573
rect 34517 25395 34518 25573
rect 34338 25394 34518 25395
rect 38338 25573 38518 25574
rect 38338 25395 38339 25573
rect 38517 25395 38518 25573
rect 38338 25394 38518 25395
rect 400 24999 580 25000
rect 400 24821 401 24999
rect 579 24821 580 24999
rect 3734 24996 3740 25002
rect 3780 24996 3786 25002
rect 4400 24999 4580 25000
rect 3728 24990 3734 24996
rect 3786 24990 3792 24996
rect 3728 24944 3734 24950
rect 3786 24944 3792 24950
rect 3734 24938 3740 24944
rect 3780 24938 3786 24944
rect 400 24820 580 24821
rect 4400 24821 4401 24999
rect 4579 24821 4580 24999
rect 7734 24996 7740 25002
rect 7780 24996 7786 25002
rect 8400 24999 8580 25000
rect 7728 24990 7734 24996
rect 7786 24990 7792 24996
rect 7728 24944 7734 24950
rect 7786 24944 7792 24950
rect 7734 24938 7740 24944
rect 7780 24938 7786 24944
rect 4400 24820 4580 24821
rect 8400 24821 8401 24999
rect 8579 24821 8580 24999
rect 11734 24996 11740 25002
rect 11780 24996 11786 25002
rect 12400 24999 12580 25000
rect 11728 24990 11734 24996
rect 11786 24990 11792 24996
rect 11728 24944 11734 24950
rect 11786 24944 11792 24950
rect 11734 24938 11740 24944
rect 11780 24938 11786 24944
rect 8400 24820 8580 24821
rect 12400 24821 12401 24999
rect 12579 24821 12580 24999
rect 15734 24996 15740 25002
rect 15780 24996 15786 25002
rect 16400 24999 16580 25000
rect 15728 24990 15734 24996
rect 15786 24990 15792 24996
rect 15728 24944 15734 24950
rect 15786 24944 15792 24950
rect 15734 24938 15740 24944
rect 15780 24938 15786 24944
rect 12400 24820 12580 24821
rect 16400 24821 16401 24999
rect 16579 24821 16580 24999
rect 19734 24996 19740 25002
rect 19780 24996 19786 25002
rect 20400 24999 20580 25000
rect 19728 24990 19734 24996
rect 19786 24990 19792 24996
rect 19728 24944 19734 24950
rect 19786 24944 19792 24950
rect 19734 24938 19740 24944
rect 19780 24938 19786 24944
rect 16400 24820 16580 24821
rect 20400 24821 20401 24999
rect 20579 24821 20580 24999
rect 23734 24996 23740 25002
rect 23780 24996 23786 25002
rect 24400 24999 24580 25000
rect 23728 24990 23734 24996
rect 23786 24990 23792 24996
rect 23728 24944 23734 24950
rect 23786 24944 23792 24950
rect 23734 24938 23740 24944
rect 23780 24938 23786 24944
rect 20400 24820 20580 24821
rect 24400 24821 24401 24999
rect 24579 24821 24580 24999
rect 27734 24996 27740 25002
rect 27780 24996 27786 25002
rect 28400 24999 28580 25000
rect 27728 24990 27734 24996
rect 27786 24990 27792 24996
rect 27728 24944 27734 24950
rect 27786 24944 27792 24950
rect 27734 24938 27740 24944
rect 27780 24938 27786 24944
rect 24400 24820 24580 24821
rect 28400 24821 28401 24999
rect 28579 24821 28580 24999
rect 31734 24996 31740 25002
rect 31780 24996 31786 25002
rect 32400 24999 32580 25000
rect 31728 24990 31734 24996
rect 31786 24990 31792 24996
rect 31728 24944 31734 24950
rect 31786 24944 31792 24950
rect 31734 24938 31740 24944
rect 31780 24938 31786 24944
rect 28400 24820 28580 24821
rect 32400 24821 32401 24999
rect 32579 24821 32580 24999
rect 35734 24996 35740 25002
rect 35780 24996 35786 25002
rect 36400 24999 36580 25000
rect 35728 24990 35734 24996
rect 35786 24990 35792 24996
rect 35728 24944 35734 24950
rect 35786 24944 35792 24950
rect 35734 24938 35740 24944
rect 35780 24938 35786 24944
rect 32400 24820 32580 24821
rect 36400 24821 36401 24999
rect 36579 24821 36580 24999
rect 39734 24996 39740 25002
rect 39780 24996 39786 25002
rect 39728 24990 39734 24996
rect 39786 24990 39792 24996
rect 39728 24944 39734 24950
rect 39786 24944 39792 24950
rect 39734 24938 39740 24944
rect 39780 24938 39786 24944
rect 36400 24820 36580 24821
rect 3262 24808 3268 24814
rect 3308 24808 3314 24814
rect 7262 24808 7268 24814
rect 7308 24808 7314 24814
rect 11262 24808 11268 24814
rect 11308 24808 11314 24814
rect 15262 24808 15268 24814
rect 15308 24808 15314 24814
rect 19262 24808 19268 24814
rect 19308 24808 19314 24814
rect 23262 24808 23268 24814
rect 23308 24808 23314 24814
rect 27262 24808 27268 24814
rect 27308 24808 27314 24814
rect 31262 24808 31268 24814
rect 31308 24808 31314 24814
rect 35262 24808 35268 24814
rect 35308 24808 35314 24814
rect 39262 24808 39268 24814
rect 39308 24808 39314 24814
rect 3256 24802 3262 24808
rect 3314 24802 3320 24808
rect 7256 24802 7262 24808
rect 7314 24802 7320 24808
rect 11256 24802 11262 24808
rect 11314 24802 11320 24808
rect 15256 24802 15262 24808
rect 15314 24802 15320 24808
rect 19256 24802 19262 24808
rect 19314 24802 19320 24808
rect 23256 24802 23262 24808
rect 23314 24802 23320 24808
rect 27256 24802 27262 24808
rect 27314 24802 27320 24808
rect 31256 24802 31262 24808
rect 31314 24802 31320 24808
rect 35256 24802 35262 24808
rect 35314 24802 35320 24808
rect 39256 24802 39262 24808
rect 39314 24802 39320 24808
rect 3256 24756 3262 24762
rect 3314 24756 3320 24762
rect 7256 24756 7262 24762
rect 7314 24756 7320 24762
rect 11256 24756 11262 24762
rect 11314 24756 11320 24762
rect 15256 24756 15262 24762
rect 15314 24756 15320 24762
rect 19256 24756 19262 24762
rect 19314 24756 19320 24762
rect 23256 24756 23262 24762
rect 23314 24756 23320 24762
rect 27256 24756 27262 24762
rect 27314 24756 27320 24762
rect 31256 24756 31262 24762
rect 31314 24756 31320 24762
rect 35256 24756 35262 24762
rect 35314 24756 35320 24762
rect 39256 24756 39262 24762
rect 39314 24756 39320 24762
rect 3262 24750 3268 24756
rect 3308 24750 3314 24756
rect 7262 24750 7268 24756
rect 7308 24750 7314 24756
rect 11262 24750 11268 24756
rect 11308 24750 11314 24756
rect 15262 24750 15268 24756
rect 15308 24750 15314 24756
rect 19262 24750 19268 24756
rect 19308 24750 19314 24756
rect 23262 24750 23268 24756
rect 23308 24750 23314 24756
rect 27262 24750 27268 24756
rect 27308 24750 27314 24756
rect 31262 24750 31268 24756
rect 31308 24750 31314 24756
rect 35262 24750 35268 24756
rect 35308 24750 35314 24756
rect 39262 24750 39268 24756
rect 39308 24750 39314 24756
rect 2240 24296 2480 24320
rect 2240 24104 2264 24296
rect 2456 24104 2480 24296
rect 2240 24080 2480 24104
rect 6240 24296 6480 24320
rect 6240 24104 6264 24296
rect 6456 24104 6480 24296
rect 6240 24080 6480 24104
rect 10240 24296 10480 24320
rect 10240 24104 10264 24296
rect 10456 24104 10480 24296
rect 10240 24080 10480 24104
rect 14240 24296 14480 24320
rect 14240 24104 14264 24296
rect 14456 24104 14480 24296
rect 14240 24080 14480 24104
rect 18240 24296 18480 24320
rect 18240 24104 18264 24296
rect 18456 24104 18480 24296
rect 18240 24080 18480 24104
rect 22240 24296 22480 24320
rect 22240 24104 22264 24296
rect 22456 24104 22480 24296
rect 22240 24080 22480 24104
rect 26240 24296 26480 24320
rect 26240 24104 26264 24296
rect 26456 24104 26480 24296
rect 26240 24080 26480 24104
rect 30240 24296 30480 24320
rect 30240 24104 30264 24296
rect 30456 24104 30480 24296
rect 30240 24080 30480 24104
rect 34240 24296 34480 24320
rect 34240 24104 34264 24296
rect 34456 24104 34480 24296
rect 34240 24080 34480 24104
rect 38240 24296 38480 24320
rect 38240 24104 38264 24296
rect 38456 24104 38480 24296
rect 38240 24080 38480 24104
rect 2240 23596 2480 23620
rect 2240 23536 2264 23596
rect 2456 23536 2480 23596
rect 2240 23380 2480 23536
rect 6240 23596 6480 23620
rect 6240 23536 6264 23596
rect 6456 23536 6480 23596
rect 6240 23380 6480 23536
rect 10240 23596 10480 23620
rect 10240 23536 10264 23596
rect 10456 23536 10480 23596
rect 10240 23380 10480 23536
rect 14240 23596 14480 23620
rect 14240 23536 14264 23596
rect 14456 23536 14480 23596
rect 14240 23380 14480 23536
rect 18240 23596 18480 23620
rect 18240 23536 18264 23596
rect 18456 23536 18480 23596
rect 18240 23380 18480 23536
rect 22240 23596 22480 23620
rect 22240 23536 22264 23596
rect 22456 23536 22480 23596
rect 22240 23380 22480 23536
rect 26240 23596 26480 23620
rect 26240 23536 26264 23596
rect 26456 23536 26480 23596
rect 26240 23380 26480 23536
rect 30240 23596 30480 23620
rect 30240 23536 30264 23596
rect 30456 23536 30480 23596
rect 30240 23380 30480 23536
rect 34240 23596 34480 23620
rect 34240 23536 34264 23596
rect 34456 23536 34480 23596
rect 34240 23380 34480 23536
rect 38240 23596 38480 23620
rect 38240 23536 38264 23596
rect 38456 23536 38480 23596
rect 38240 23380 38480 23536
rect 1936 23160 2256 23216
rect 360 22916 600 22940
rect 360 22724 384 22916
rect 576 22724 600 22916
rect 1936 22920 1960 23160
rect 2224 22920 2256 23160
rect 3602 23163 3690 23168
rect 3602 23085 3607 23163
rect 3685 23085 3690 23163
rect 3602 23080 3690 23085
rect 5936 23160 6256 23216
rect 1936 22896 2256 22920
rect 4360 22916 4600 22940
rect 360 22700 600 22724
rect 4360 22724 4384 22916
rect 4576 22724 4600 22916
rect 5936 22920 5960 23160
rect 6224 22920 6256 23160
rect 7602 23163 7690 23168
rect 7602 23085 7607 23163
rect 7685 23085 7690 23163
rect 7602 23080 7690 23085
rect 9936 23160 10256 23216
rect 5936 22896 6256 22920
rect 8360 22916 8600 22940
rect 2810 22711 2946 22716
rect 2810 22637 2815 22711
rect 2941 22637 2946 22711
rect 4360 22700 4600 22724
rect 8360 22724 8384 22916
rect 8576 22724 8600 22916
rect 9936 22920 9960 23160
rect 10224 22920 10256 23160
rect 11602 23163 11690 23168
rect 11602 23085 11607 23163
rect 11685 23085 11690 23163
rect 11602 23080 11690 23085
rect 13936 23160 14256 23216
rect 9936 22896 10256 22920
rect 12360 22916 12600 22940
rect 6810 22711 6946 22716
rect 2810 22632 2946 22637
rect 6810 22637 6815 22711
rect 6941 22637 6946 22711
rect 8360 22700 8600 22724
rect 12360 22724 12384 22916
rect 12576 22724 12600 22916
rect 13936 22920 13960 23160
rect 14224 22920 14256 23160
rect 15602 23163 15690 23168
rect 15602 23085 15607 23163
rect 15685 23085 15690 23163
rect 15602 23080 15690 23085
rect 17936 23160 18256 23216
rect 13936 22896 14256 22920
rect 16360 22916 16600 22940
rect 10810 22711 10946 22716
rect 6810 22632 6946 22637
rect 10810 22637 10815 22711
rect 10941 22637 10946 22711
rect 12360 22700 12600 22724
rect 16360 22724 16384 22916
rect 16576 22724 16600 22916
rect 17936 22920 17960 23160
rect 18224 22920 18256 23160
rect 19602 23163 19690 23168
rect 19602 23085 19607 23163
rect 19685 23085 19690 23163
rect 19602 23080 19690 23085
rect 21936 23160 22256 23216
rect 17936 22896 18256 22920
rect 20360 22916 20600 22940
rect 14810 22711 14946 22716
rect 10810 22632 10946 22637
rect 14810 22637 14815 22711
rect 14941 22637 14946 22711
rect 16360 22700 16600 22724
rect 20360 22724 20384 22916
rect 20576 22724 20600 22916
rect 21936 22920 21960 23160
rect 22224 22920 22256 23160
rect 23602 23163 23690 23168
rect 23602 23085 23607 23163
rect 23685 23085 23690 23163
rect 23602 23080 23690 23085
rect 25936 23160 26256 23216
rect 21936 22896 22256 22920
rect 24360 22916 24600 22940
rect 18810 22711 18946 22716
rect 14810 22632 14946 22637
rect 18810 22637 18815 22711
rect 18941 22637 18946 22711
rect 20360 22700 20600 22724
rect 24360 22724 24384 22916
rect 24576 22724 24600 22916
rect 25936 22920 25960 23160
rect 26224 22920 26256 23160
rect 27602 23163 27690 23168
rect 27602 23085 27607 23163
rect 27685 23085 27690 23163
rect 27602 23080 27690 23085
rect 29936 23160 30256 23216
rect 25936 22896 26256 22920
rect 28360 22916 28600 22940
rect 22810 22711 22946 22716
rect 18810 22632 18946 22637
rect 22810 22637 22815 22711
rect 22941 22637 22946 22711
rect 24360 22700 24600 22724
rect 28360 22724 28384 22916
rect 28576 22724 28600 22916
rect 29936 22920 29960 23160
rect 30224 22920 30256 23160
rect 31602 23163 31690 23168
rect 31602 23085 31607 23163
rect 31685 23085 31690 23163
rect 31602 23080 31690 23085
rect 33936 23160 34256 23216
rect 29936 22896 30256 22920
rect 32360 22916 32600 22940
rect 26810 22711 26946 22716
rect 22810 22632 22946 22637
rect 26810 22637 26815 22711
rect 26941 22637 26946 22711
rect 28360 22700 28600 22724
rect 32360 22724 32384 22916
rect 32576 22724 32600 22916
rect 33936 22920 33960 23160
rect 34224 22920 34256 23160
rect 35602 23163 35690 23168
rect 35602 23085 35607 23163
rect 35685 23085 35690 23163
rect 35602 23080 35690 23085
rect 37936 23160 38256 23216
rect 33936 22896 34256 22920
rect 36360 22916 36600 22940
rect 30810 22711 30946 22716
rect 26810 22632 26946 22637
rect 30810 22637 30815 22711
rect 30941 22637 30946 22711
rect 32360 22700 32600 22724
rect 36360 22724 36384 22916
rect 36576 22724 36600 22916
rect 37936 22920 37960 23160
rect 38224 22920 38256 23160
rect 39602 23163 39690 23168
rect 39602 23085 39607 23163
rect 39685 23085 39690 23163
rect 39602 23080 39690 23085
rect 37936 22896 38256 22920
rect 34810 22711 34946 22716
rect 30810 22632 30946 22637
rect 34810 22637 34815 22711
rect 34941 22637 34946 22711
rect 36360 22700 36600 22724
rect 38810 22711 38946 22716
rect 34810 22632 34946 22637
rect 38810 22637 38815 22711
rect 38941 22637 38946 22711
rect 38810 22632 38946 22637
rect 2338 22573 2518 22574
rect 2338 22395 2339 22573
rect 2517 22395 2518 22573
rect 2338 22394 2518 22395
rect 6338 22573 6518 22574
rect 6338 22395 6339 22573
rect 6517 22395 6518 22573
rect 6338 22394 6518 22395
rect 10338 22573 10518 22574
rect 10338 22395 10339 22573
rect 10517 22395 10518 22573
rect 10338 22394 10518 22395
rect 14338 22573 14518 22574
rect 14338 22395 14339 22573
rect 14517 22395 14518 22573
rect 14338 22394 14518 22395
rect 18338 22573 18518 22574
rect 18338 22395 18339 22573
rect 18517 22395 18518 22573
rect 18338 22394 18518 22395
rect 22338 22573 22518 22574
rect 22338 22395 22339 22573
rect 22517 22395 22518 22573
rect 22338 22394 22518 22395
rect 26338 22573 26518 22574
rect 26338 22395 26339 22573
rect 26517 22395 26518 22573
rect 26338 22394 26518 22395
rect 30338 22573 30518 22574
rect 30338 22395 30339 22573
rect 30517 22395 30518 22573
rect 30338 22394 30518 22395
rect 34338 22573 34518 22574
rect 34338 22395 34339 22573
rect 34517 22395 34518 22573
rect 34338 22394 34518 22395
rect 38338 22573 38518 22574
rect 38338 22395 38339 22573
rect 38517 22395 38518 22573
rect 38338 22394 38518 22395
rect 400 21999 580 22000
rect 400 21821 401 21999
rect 579 21821 580 21999
rect 3734 21996 3740 22002
rect 3780 21996 3786 22002
rect 4400 21999 4580 22000
rect 3728 21990 3734 21996
rect 3786 21990 3792 21996
rect 3728 21944 3734 21950
rect 3786 21944 3792 21950
rect 3734 21938 3740 21944
rect 3780 21938 3786 21944
rect 400 21820 580 21821
rect 4400 21821 4401 21999
rect 4579 21821 4580 21999
rect 7734 21996 7740 22002
rect 7780 21996 7786 22002
rect 8400 21999 8580 22000
rect 7728 21990 7734 21996
rect 7786 21990 7792 21996
rect 7728 21944 7734 21950
rect 7786 21944 7792 21950
rect 7734 21938 7740 21944
rect 7780 21938 7786 21944
rect 4400 21820 4580 21821
rect 8400 21821 8401 21999
rect 8579 21821 8580 21999
rect 11734 21996 11740 22002
rect 11780 21996 11786 22002
rect 12400 21999 12580 22000
rect 11728 21990 11734 21996
rect 11786 21990 11792 21996
rect 11728 21944 11734 21950
rect 11786 21944 11792 21950
rect 11734 21938 11740 21944
rect 11780 21938 11786 21944
rect 8400 21820 8580 21821
rect 12400 21821 12401 21999
rect 12579 21821 12580 21999
rect 15734 21996 15740 22002
rect 15780 21996 15786 22002
rect 16400 21999 16580 22000
rect 15728 21990 15734 21996
rect 15786 21990 15792 21996
rect 15728 21944 15734 21950
rect 15786 21944 15792 21950
rect 15734 21938 15740 21944
rect 15780 21938 15786 21944
rect 12400 21820 12580 21821
rect 16400 21821 16401 21999
rect 16579 21821 16580 21999
rect 19734 21996 19740 22002
rect 19780 21996 19786 22002
rect 20400 21999 20580 22000
rect 19728 21990 19734 21996
rect 19786 21990 19792 21996
rect 19728 21944 19734 21950
rect 19786 21944 19792 21950
rect 19734 21938 19740 21944
rect 19780 21938 19786 21944
rect 16400 21820 16580 21821
rect 20400 21821 20401 21999
rect 20579 21821 20580 21999
rect 23734 21996 23740 22002
rect 23780 21996 23786 22002
rect 24400 21999 24580 22000
rect 23728 21990 23734 21996
rect 23786 21990 23792 21996
rect 23728 21944 23734 21950
rect 23786 21944 23792 21950
rect 23734 21938 23740 21944
rect 23780 21938 23786 21944
rect 20400 21820 20580 21821
rect 24400 21821 24401 21999
rect 24579 21821 24580 21999
rect 27734 21996 27740 22002
rect 27780 21996 27786 22002
rect 28400 21999 28580 22000
rect 27728 21990 27734 21996
rect 27786 21990 27792 21996
rect 27728 21944 27734 21950
rect 27786 21944 27792 21950
rect 27734 21938 27740 21944
rect 27780 21938 27786 21944
rect 24400 21820 24580 21821
rect 28400 21821 28401 21999
rect 28579 21821 28580 21999
rect 31734 21996 31740 22002
rect 31780 21996 31786 22002
rect 32400 21999 32580 22000
rect 31728 21990 31734 21996
rect 31786 21990 31792 21996
rect 31728 21944 31734 21950
rect 31786 21944 31792 21950
rect 31734 21938 31740 21944
rect 31780 21938 31786 21944
rect 28400 21820 28580 21821
rect 32400 21821 32401 21999
rect 32579 21821 32580 21999
rect 35734 21996 35740 22002
rect 35780 21996 35786 22002
rect 36400 21999 36580 22000
rect 35728 21990 35734 21996
rect 35786 21990 35792 21996
rect 35728 21944 35734 21950
rect 35786 21944 35792 21950
rect 35734 21938 35740 21944
rect 35780 21938 35786 21944
rect 32400 21820 32580 21821
rect 36400 21821 36401 21999
rect 36579 21821 36580 21999
rect 39734 21996 39740 22002
rect 39780 21996 39786 22002
rect 39728 21990 39734 21996
rect 39786 21990 39792 21996
rect 39728 21944 39734 21950
rect 39786 21944 39792 21950
rect 39734 21938 39740 21944
rect 39780 21938 39786 21944
rect 36400 21820 36580 21821
rect 3262 21808 3268 21814
rect 3308 21808 3314 21814
rect 7262 21808 7268 21814
rect 7308 21808 7314 21814
rect 11262 21808 11268 21814
rect 11308 21808 11314 21814
rect 15262 21808 15268 21814
rect 15308 21808 15314 21814
rect 19262 21808 19268 21814
rect 19308 21808 19314 21814
rect 23262 21808 23268 21814
rect 23308 21808 23314 21814
rect 27262 21808 27268 21814
rect 27308 21808 27314 21814
rect 31262 21808 31268 21814
rect 31308 21808 31314 21814
rect 35262 21808 35268 21814
rect 35308 21808 35314 21814
rect 39262 21808 39268 21814
rect 39308 21808 39314 21814
rect 3256 21802 3262 21808
rect 3314 21802 3320 21808
rect 7256 21802 7262 21808
rect 7314 21802 7320 21808
rect 11256 21802 11262 21808
rect 11314 21802 11320 21808
rect 15256 21802 15262 21808
rect 15314 21802 15320 21808
rect 19256 21802 19262 21808
rect 19314 21802 19320 21808
rect 23256 21802 23262 21808
rect 23314 21802 23320 21808
rect 27256 21802 27262 21808
rect 27314 21802 27320 21808
rect 31256 21802 31262 21808
rect 31314 21802 31320 21808
rect 35256 21802 35262 21808
rect 35314 21802 35320 21808
rect 39256 21802 39262 21808
rect 39314 21802 39320 21808
rect 3256 21756 3262 21762
rect 3314 21756 3320 21762
rect 7256 21756 7262 21762
rect 7314 21756 7320 21762
rect 11256 21756 11262 21762
rect 11314 21756 11320 21762
rect 15256 21756 15262 21762
rect 15314 21756 15320 21762
rect 19256 21756 19262 21762
rect 19314 21756 19320 21762
rect 23256 21756 23262 21762
rect 23314 21756 23320 21762
rect 27256 21756 27262 21762
rect 27314 21756 27320 21762
rect 31256 21756 31262 21762
rect 31314 21756 31320 21762
rect 35256 21756 35262 21762
rect 35314 21756 35320 21762
rect 39256 21756 39262 21762
rect 39314 21756 39320 21762
rect 3262 21750 3268 21756
rect 3308 21750 3314 21756
rect 7262 21750 7268 21756
rect 7308 21750 7314 21756
rect 11262 21750 11268 21756
rect 11308 21750 11314 21756
rect 15262 21750 15268 21756
rect 15308 21750 15314 21756
rect 19262 21750 19268 21756
rect 19308 21750 19314 21756
rect 23262 21750 23268 21756
rect 23308 21750 23314 21756
rect 27262 21750 27268 21756
rect 27308 21750 27314 21756
rect 31262 21750 31268 21756
rect 31308 21750 31314 21756
rect 35262 21750 35268 21756
rect 35308 21750 35314 21756
rect 39262 21750 39268 21756
rect 39308 21750 39314 21756
rect 2240 21296 2480 21320
rect 2240 21104 2264 21296
rect 2456 21104 2480 21296
rect 2240 21080 2480 21104
rect 6240 21296 6480 21320
rect 6240 21104 6264 21296
rect 6456 21104 6480 21296
rect 6240 21080 6480 21104
rect 10240 21296 10480 21320
rect 10240 21104 10264 21296
rect 10456 21104 10480 21296
rect 10240 21080 10480 21104
rect 14240 21296 14480 21320
rect 14240 21104 14264 21296
rect 14456 21104 14480 21296
rect 14240 21080 14480 21104
rect 18240 21296 18480 21320
rect 18240 21104 18264 21296
rect 18456 21104 18480 21296
rect 18240 21080 18480 21104
rect 22240 21296 22480 21320
rect 22240 21104 22264 21296
rect 22456 21104 22480 21296
rect 22240 21080 22480 21104
rect 26240 21296 26480 21320
rect 26240 21104 26264 21296
rect 26456 21104 26480 21296
rect 26240 21080 26480 21104
rect 30240 21296 30480 21320
rect 30240 21104 30264 21296
rect 30456 21104 30480 21296
rect 30240 21080 30480 21104
rect 34240 21296 34480 21320
rect 34240 21104 34264 21296
rect 34456 21104 34480 21296
rect 34240 21080 34480 21104
rect 38240 21296 38480 21320
rect 38240 21104 38264 21296
rect 38456 21104 38480 21296
rect 38240 21080 38480 21104
rect 2240 20596 2480 20620
rect 2240 20536 2264 20596
rect 2456 20536 2480 20596
rect 2240 20380 2480 20536
rect 6240 20596 6480 20620
rect 6240 20536 6264 20596
rect 6456 20536 6480 20596
rect 6240 20380 6480 20536
rect 10240 20596 10480 20620
rect 10240 20536 10264 20596
rect 10456 20536 10480 20596
rect 10240 20380 10480 20536
rect 14240 20596 14480 20620
rect 14240 20536 14264 20596
rect 14456 20536 14480 20596
rect 14240 20380 14480 20536
rect 18240 20596 18480 20620
rect 18240 20536 18264 20596
rect 18456 20536 18480 20596
rect 18240 20380 18480 20536
rect 22240 20596 22480 20620
rect 22240 20536 22264 20596
rect 22456 20536 22480 20596
rect 22240 20380 22480 20536
rect 26240 20596 26480 20620
rect 26240 20536 26264 20596
rect 26456 20536 26480 20596
rect 26240 20380 26480 20536
rect 30240 20596 30480 20620
rect 30240 20536 30264 20596
rect 30456 20536 30480 20596
rect 30240 20380 30480 20536
rect 34240 20596 34480 20620
rect 34240 20536 34264 20596
rect 34456 20536 34480 20596
rect 34240 20380 34480 20536
rect 38240 20596 38480 20620
rect 38240 20536 38264 20596
rect 38456 20536 38480 20596
rect 38240 20380 38480 20536
rect 1936 20160 2256 20216
rect 360 19916 600 19940
rect 360 19724 384 19916
rect 576 19724 600 19916
rect 1936 19920 1960 20160
rect 2224 19920 2256 20160
rect 3602 20163 3690 20168
rect 3602 20085 3607 20163
rect 3685 20085 3690 20163
rect 3602 20080 3690 20085
rect 5936 20160 6256 20216
rect 1936 19896 2256 19920
rect 4360 19916 4600 19940
rect 360 19700 600 19724
rect 4360 19724 4384 19916
rect 4576 19724 4600 19916
rect 5936 19920 5960 20160
rect 6224 19920 6256 20160
rect 7602 20163 7690 20168
rect 7602 20085 7607 20163
rect 7685 20085 7690 20163
rect 7602 20080 7690 20085
rect 9936 20160 10256 20216
rect 5936 19896 6256 19920
rect 8360 19916 8600 19940
rect 2810 19711 2946 19716
rect 2810 19637 2815 19711
rect 2941 19637 2946 19711
rect 4360 19700 4600 19724
rect 8360 19724 8384 19916
rect 8576 19724 8600 19916
rect 9936 19920 9960 20160
rect 10224 19920 10256 20160
rect 11602 20163 11690 20168
rect 11602 20085 11607 20163
rect 11685 20085 11690 20163
rect 11602 20080 11690 20085
rect 13936 20160 14256 20216
rect 9936 19896 10256 19920
rect 12360 19916 12600 19940
rect 6810 19711 6946 19716
rect 2810 19632 2946 19637
rect 6810 19637 6815 19711
rect 6941 19637 6946 19711
rect 8360 19700 8600 19724
rect 12360 19724 12384 19916
rect 12576 19724 12600 19916
rect 13936 19920 13960 20160
rect 14224 19920 14256 20160
rect 15602 20163 15690 20168
rect 15602 20085 15607 20163
rect 15685 20085 15690 20163
rect 15602 20080 15690 20085
rect 17936 20160 18256 20216
rect 13936 19896 14256 19920
rect 16360 19916 16600 19940
rect 10810 19711 10946 19716
rect 6810 19632 6946 19637
rect 10810 19637 10815 19711
rect 10941 19637 10946 19711
rect 12360 19700 12600 19724
rect 16360 19724 16384 19916
rect 16576 19724 16600 19916
rect 17936 19920 17960 20160
rect 18224 19920 18256 20160
rect 19602 20163 19690 20168
rect 19602 20085 19607 20163
rect 19685 20085 19690 20163
rect 19602 20080 19690 20085
rect 21936 20160 22256 20216
rect 17936 19896 18256 19920
rect 20360 19916 20600 19940
rect 14810 19711 14946 19716
rect 10810 19632 10946 19637
rect 14810 19637 14815 19711
rect 14941 19637 14946 19711
rect 16360 19700 16600 19724
rect 20360 19724 20384 19916
rect 20576 19724 20600 19916
rect 21936 19920 21960 20160
rect 22224 19920 22256 20160
rect 23602 20163 23690 20168
rect 23602 20085 23607 20163
rect 23685 20085 23690 20163
rect 23602 20080 23690 20085
rect 25936 20160 26256 20216
rect 21936 19896 22256 19920
rect 24360 19916 24600 19940
rect 18810 19711 18946 19716
rect 14810 19632 14946 19637
rect 18810 19637 18815 19711
rect 18941 19637 18946 19711
rect 20360 19700 20600 19724
rect 24360 19724 24384 19916
rect 24576 19724 24600 19916
rect 25936 19920 25960 20160
rect 26224 19920 26256 20160
rect 27602 20163 27690 20168
rect 27602 20085 27607 20163
rect 27685 20085 27690 20163
rect 27602 20080 27690 20085
rect 29936 20160 30256 20216
rect 25936 19896 26256 19920
rect 28360 19916 28600 19940
rect 22810 19711 22946 19716
rect 18810 19632 18946 19637
rect 22810 19637 22815 19711
rect 22941 19637 22946 19711
rect 24360 19700 24600 19724
rect 28360 19724 28384 19916
rect 28576 19724 28600 19916
rect 29936 19920 29960 20160
rect 30224 19920 30256 20160
rect 31602 20163 31690 20168
rect 31602 20085 31607 20163
rect 31685 20085 31690 20163
rect 31602 20080 31690 20085
rect 33936 20160 34256 20216
rect 29936 19896 30256 19920
rect 32360 19916 32600 19940
rect 26810 19711 26946 19716
rect 22810 19632 22946 19637
rect 26810 19637 26815 19711
rect 26941 19637 26946 19711
rect 28360 19700 28600 19724
rect 32360 19724 32384 19916
rect 32576 19724 32600 19916
rect 33936 19920 33960 20160
rect 34224 19920 34256 20160
rect 35602 20163 35690 20168
rect 35602 20085 35607 20163
rect 35685 20085 35690 20163
rect 35602 20080 35690 20085
rect 37936 20160 38256 20216
rect 33936 19896 34256 19920
rect 36360 19916 36600 19940
rect 30810 19711 30946 19716
rect 26810 19632 26946 19637
rect 30810 19637 30815 19711
rect 30941 19637 30946 19711
rect 32360 19700 32600 19724
rect 36360 19724 36384 19916
rect 36576 19724 36600 19916
rect 37936 19920 37960 20160
rect 38224 19920 38256 20160
rect 39602 20163 39690 20168
rect 39602 20085 39607 20163
rect 39685 20085 39690 20163
rect 39602 20080 39690 20085
rect 37936 19896 38256 19920
rect 34810 19711 34946 19716
rect 30810 19632 30946 19637
rect 34810 19637 34815 19711
rect 34941 19637 34946 19711
rect 36360 19700 36600 19724
rect 38810 19711 38946 19716
rect 34810 19632 34946 19637
rect 38810 19637 38815 19711
rect 38941 19637 38946 19711
rect 38810 19632 38946 19637
rect 2338 19573 2518 19574
rect 2338 19395 2339 19573
rect 2517 19395 2518 19573
rect 2338 19394 2518 19395
rect 6338 19573 6518 19574
rect 6338 19395 6339 19573
rect 6517 19395 6518 19573
rect 6338 19394 6518 19395
rect 10338 19573 10518 19574
rect 10338 19395 10339 19573
rect 10517 19395 10518 19573
rect 10338 19394 10518 19395
rect 14338 19573 14518 19574
rect 14338 19395 14339 19573
rect 14517 19395 14518 19573
rect 14338 19394 14518 19395
rect 18338 19573 18518 19574
rect 18338 19395 18339 19573
rect 18517 19395 18518 19573
rect 18338 19394 18518 19395
rect 22338 19573 22518 19574
rect 22338 19395 22339 19573
rect 22517 19395 22518 19573
rect 22338 19394 22518 19395
rect 26338 19573 26518 19574
rect 26338 19395 26339 19573
rect 26517 19395 26518 19573
rect 26338 19394 26518 19395
rect 30338 19573 30518 19574
rect 30338 19395 30339 19573
rect 30517 19395 30518 19573
rect 30338 19394 30518 19395
rect 34338 19573 34518 19574
rect 34338 19395 34339 19573
rect 34517 19395 34518 19573
rect 34338 19394 34518 19395
rect 38338 19573 38518 19574
rect 38338 19395 38339 19573
rect 38517 19395 38518 19573
rect 38338 19394 38518 19395
rect 400 18999 580 19000
rect 400 18821 401 18999
rect 579 18821 580 18999
rect 3734 18996 3740 19002
rect 3780 18996 3786 19002
rect 4400 18999 4580 19000
rect 3728 18990 3734 18996
rect 3786 18990 3792 18996
rect 3728 18944 3734 18950
rect 3786 18944 3792 18950
rect 3734 18938 3740 18944
rect 3780 18938 3786 18944
rect 400 18820 580 18821
rect 4400 18821 4401 18999
rect 4579 18821 4580 18999
rect 7734 18996 7740 19002
rect 7780 18996 7786 19002
rect 8400 18999 8580 19000
rect 7728 18990 7734 18996
rect 7786 18990 7792 18996
rect 7728 18944 7734 18950
rect 7786 18944 7792 18950
rect 7734 18938 7740 18944
rect 7780 18938 7786 18944
rect 4400 18820 4580 18821
rect 8400 18821 8401 18999
rect 8579 18821 8580 18999
rect 11734 18996 11740 19002
rect 11780 18996 11786 19002
rect 12400 18999 12580 19000
rect 11728 18990 11734 18996
rect 11786 18990 11792 18996
rect 11728 18944 11734 18950
rect 11786 18944 11792 18950
rect 11734 18938 11740 18944
rect 11780 18938 11786 18944
rect 8400 18820 8580 18821
rect 12400 18821 12401 18999
rect 12579 18821 12580 18999
rect 15734 18996 15740 19002
rect 15780 18996 15786 19002
rect 16400 18999 16580 19000
rect 15728 18990 15734 18996
rect 15786 18990 15792 18996
rect 15728 18944 15734 18950
rect 15786 18944 15792 18950
rect 15734 18938 15740 18944
rect 15780 18938 15786 18944
rect 12400 18820 12580 18821
rect 16400 18821 16401 18999
rect 16579 18821 16580 18999
rect 19734 18996 19740 19002
rect 19780 18996 19786 19002
rect 20400 18999 20580 19000
rect 19728 18990 19734 18996
rect 19786 18990 19792 18996
rect 19728 18944 19734 18950
rect 19786 18944 19792 18950
rect 19734 18938 19740 18944
rect 19780 18938 19786 18944
rect 16400 18820 16580 18821
rect 20400 18821 20401 18999
rect 20579 18821 20580 18999
rect 23734 18996 23740 19002
rect 23780 18996 23786 19002
rect 24400 18999 24580 19000
rect 23728 18990 23734 18996
rect 23786 18990 23792 18996
rect 23728 18944 23734 18950
rect 23786 18944 23792 18950
rect 23734 18938 23740 18944
rect 23780 18938 23786 18944
rect 20400 18820 20580 18821
rect 24400 18821 24401 18999
rect 24579 18821 24580 18999
rect 27734 18996 27740 19002
rect 27780 18996 27786 19002
rect 28400 18999 28580 19000
rect 27728 18990 27734 18996
rect 27786 18990 27792 18996
rect 27728 18944 27734 18950
rect 27786 18944 27792 18950
rect 27734 18938 27740 18944
rect 27780 18938 27786 18944
rect 24400 18820 24580 18821
rect 28400 18821 28401 18999
rect 28579 18821 28580 18999
rect 31734 18996 31740 19002
rect 31780 18996 31786 19002
rect 32400 18999 32580 19000
rect 31728 18990 31734 18996
rect 31786 18990 31792 18996
rect 31728 18944 31734 18950
rect 31786 18944 31792 18950
rect 31734 18938 31740 18944
rect 31780 18938 31786 18944
rect 28400 18820 28580 18821
rect 32400 18821 32401 18999
rect 32579 18821 32580 18999
rect 35734 18996 35740 19002
rect 35780 18996 35786 19002
rect 36400 18999 36580 19000
rect 35728 18990 35734 18996
rect 35786 18990 35792 18996
rect 35728 18944 35734 18950
rect 35786 18944 35792 18950
rect 35734 18938 35740 18944
rect 35780 18938 35786 18944
rect 32400 18820 32580 18821
rect 36400 18821 36401 18999
rect 36579 18821 36580 18999
rect 39734 18996 39740 19002
rect 39780 18996 39786 19002
rect 39728 18990 39734 18996
rect 39786 18990 39792 18996
rect 39728 18944 39734 18950
rect 39786 18944 39792 18950
rect 39734 18938 39740 18944
rect 39780 18938 39786 18944
rect 36400 18820 36580 18821
rect 3262 18808 3268 18814
rect 3308 18808 3314 18814
rect 7262 18808 7268 18814
rect 7308 18808 7314 18814
rect 11262 18808 11268 18814
rect 11308 18808 11314 18814
rect 15262 18808 15268 18814
rect 15308 18808 15314 18814
rect 19262 18808 19268 18814
rect 19308 18808 19314 18814
rect 23262 18808 23268 18814
rect 23308 18808 23314 18814
rect 27262 18808 27268 18814
rect 27308 18808 27314 18814
rect 31262 18808 31268 18814
rect 31308 18808 31314 18814
rect 35262 18808 35268 18814
rect 35308 18808 35314 18814
rect 39262 18808 39268 18814
rect 39308 18808 39314 18814
rect 3256 18802 3262 18808
rect 3314 18802 3320 18808
rect 7256 18802 7262 18808
rect 7314 18802 7320 18808
rect 11256 18802 11262 18808
rect 11314 18802 11320 18808
rect 15256 18802 15262 18808
rect 15314 18802 15320 18808
rect 19256 18802 19262 18808
rect 19314 18802 19320 18808
rect 23256 18802 23262 18808
rect 23314 18802 23320 18808
rect 27256 18802 27262 18808
rect 27314 18802 27320 18808
rect 31256 18802 31262 18808
rect 31314 18802 31320 18808
rect 35256 18802 35262 18808
rect 35314 18802 35320 18808
rect 39256 18802 39262 18808
rect 39314 18802 39320 18808
rect 3256 18756 3262 18762
rect 3314 18756 3320 18762
rect 7256 18756 7262 18762
rect 7314 18756 7320 18762
rect 11256 18756 11262 18762
rect 11314 18756 11320 18762
rect 15256 18756 15262 18762
rect 15314 18756 15320 18762
rect 19256 18756 19262 18762
rect 19314 18756 19320 18762
rect 23256 18756 23262 18762
rect 23314 18756 23320 18762
rect 27256 18756 27262 18762
rect 27314 18756 27320 18762
rect 31256 18756 31262 18762
rect 31314 18756 31320 18762
rect 35256 18756 35262 18762
rect 35314 18756 35320 18762
rect 39256 18756 39262 18762
rect 39314 18756 39320 18762
rect 3262 18750 3268 18756
rect 3308 18750 3314 18756
rect 7262 18750 7268 18756
rect 7308 18750 7314 18756
rect 11262 18750 11268 18756
rect 11308 18750 11314 18756
rect 15262 18750 15268 18756
rect 15308 18750 15314 18756
rect 19262 18750 19268 18756
rect 19308 18750 19314 18756
rect 23262 18750 23268 18756
rect 23308 18750 23314 18756
rect 27262 18750 27268 18756
rect 27308 18750 27314 18756
rect 31262 18750 31268 18756
rect 31308 18750 31314 18756
rect 35262 18750 35268 18756
rect 35308 18750 35314 18756
rect 39262 18750 39268 18756
rect 39308 18750 39314 18756
rect 2240 18296 2480 18320
rect 2240 18104 2264 18296
rect 2456 18104 2480 18296
rect 2240 18080 2480 18104
rect 6240 18296 6480 18320
rect 6240 18104 6264 18296
rect 6456 18104 6480 18296
rect 6240 18080 6480 18104
rect 10240 18296 10480 18320
rect 10240 18104 10264 18296
rect 10456 18104 10480 18296
rect 10240 18080 10480 18104
rect 14240 18296 14480 18320
rect 14240 18104 14264 18296
rect 14456 18104 14480 18296
rect 14240 18080 14480 18104
rect 18240 18296 18480 18320
rect 18240 18104 18264 18296
rect 18456 18104 18480 18296
rect 18240 18080 18480 18104
rect 22240 18296 22480 18320
rect 22240 18104 22264 18296
rect 22456 18104 22480 18296
rect 22240 18080 22480 18104
rect 26240 18296 26480 18320
rect 26240 18104 26264 18296
rect 26456 18104 26480 18296
rect 26240 18080 26480 18104
rect 30240 18296 30480 18320
rect 30240 18104 30264 18296
rect 30456 18104 30480 18296
rect 30240 18080 30480 18104
rect 34240 18296 34480 18320
rect 34240 18104 34264 18296
rect 34456 18104 34480 18296
rect 34240 18080 34480 18104
rect 38240 18296 38480 18320
rect 38240 18104 38264 18296
rect 38456 18104 38480 18296
rect 38240 18080 38480 18104
rect 2240 17596 2480 17620
rect 2240 17536 2264 17596
rect 2456 17536 2480 17596
rect 2240 17380 2480 17536
rect 6240 17596 6480 17620
rect 6240 17536 6264 17596
rect 6456 17536 6480 17596
rect 6240 17380 6480 17536
rect 10240 17596 10480 17620
rect 10240 17536 10264 17596
rect 10456 17536 10480 17596
rect 10240 17380 10480 17536
rect 14240 17596 14480 17620
rect 14240 17536 14264 17596
rect 14456 17536 14480 17596
rect 14240 17380 14480 17536
rect 18240 17596 18480 17620
rect 18240 17536 18264 17596
rect 18456 17536 18480 17596
rect 18240 17380 18480 17536
rect 22240 17596 22480 17620
rect 22240 17536 22264 17596
rect 22456 17536 22480 17596
rect 22240 17380 22480 17536
rect 26240 17596 26480 17620
rect 26240 17536 26264 17596
rect 26456 17536 26480 17596
rect 26240 17380 26480 17536
rect 30240 17596 30480 17620
rect 30240 17536 30264 17596
rect 30456 17536 30480 17596
rect 30240 17380 30480 17536
rect 34240 17596 34480 17620
rect 34240 17536 34264 17596
rect 34456 17536 34480 17596
rect 34240 17380 34480 17536
rect 38240 17596 38480 17620
rect 38240 17536 38264 17596
rect 38456 17536 38480 17596
rect 38240 17380 38480 17536
rect 1936 17160 2256 17216
rect 360 16916 600 16940
rect 360 16724 384 16916
rect 576 16724 600 16916
rect 1936 16920 1960 17160
rect 2224 16920 2256 17160
rect 3602 17163 3690 17168
rect 3602 17085 3607 17163
rect 3685 17085 3690 17163
rect 3602 17080 3690 17085
rect 5936 17160 6256 17216
rect 1936 16896 2256 16920
rect 4360 16916 4600 16940
rect 360 16700 600 16724
rect 4360 16724 4384 16916
rect 4576 16724 4600 16916
rect 5936 16920 5960 17160
rect 6224 16920 6256 17160
rect 7602 17163 7690 17168
rect 7602 17085 7607 17163
rect 7685 17085 7690 17163
rect 7602 17080 7690 17085
rect 9936 17160 10256 17216
rect 5936 16896 6256 16920
rect 8360 16916 8600 16940
rect 2810 16711 2946 16716
rect 2810 16637 2815 16711
rect 2941 16637 2946 16711
rect 4360 16700 4600 16724
rect 8360 16724 8384 16916
rect 8576 16724 8600 16916
rect 9936 16920 9960 17160
rect 10224 16920 10256 17160
rect 11602 17163 11690 17168
rect 11602 17085 11607 17163
rect 11685 17085 11690 17163
rect 11602 17080 11690 17085
rect 13936 17160 14256 17216
rect 9936 16896 10256 16920
rect 12360 16916 12600 16940
rect 6810 16711 6946 16716
rect 2810 16632 2946 16637
rect 6810 16637 6815 16711
rect 6941 16637 6946 16711
rect 8360 16700 8600 16724
rect 12360 16724 12384 16916
rect 12576 16724 12600 16916
rect 13936 16920 13960 17160
rect 14224 16920 14256 17160
rect 15602 17163 15690 17168
rect 15602 17085 15607 17163
rect 15685 17085 15690 17163
rect 15602 17080 15690 17085
rect 17936 17160 18256 17216
rect 13936 16896 14256 16920
rect 16360 16916 16600 16940
rect 10810 16711 10946 16716
rect 6810 16632 6946 16637
rect 10810 16637 10815 16711
rect 10941 16637 10946 16711
rect 12360 16700 12600 16724
rect 16360 16724 16384 16916
rect 16576 16724 16600 16916
rect 17936 16920 17960 17160
rect 18224 16920 18256 17160
rect 19602 17163 19690 17168
rect 19602 17085 19607 17163
rect 19685 17085 19690 17163
rect 19602 17080 19690 17085
rect 21936 17160 22256 17216
rect 17936 16896 18256 16920
rect 20360 16916 20600 16940
rect 14810 16711 14946 16716
rect 10810 16632 10946 16637
rect 14810 16637 14815 16711
rect 14941 16637 14946 16711
rect 16360 16700 16600 16724
rect 20360 16724 20384 16916
rect 20576 16724 20600 16916
rect 21936 16920 21960 17160
rect 22224 16920 22256 17160
rect 23602 17163 23690 17168
rect 23602 17085 23607 17163
rect 23685 17085 23690 17163
rect 23602 17080 23690 17085
rect 25936 17160 26256 17216
rect 21936 16896 22256 16920
rect 24360 16916 24600 16940
rect 18810 16711 18946 16716
rect 14810 16632 14946 16637
rect 18810 16637 18815 16711
rect 18941 16637 18946 16711
rect 20360 16700 20600 16724
rect 24360 16724 24384 16916
rect 24576 16724 24600 16916
rect 25936 16920 25960 17160
rect 26224 16920 26256 17160
rect 27602 17163 27690 17168
rect 27602 17085 27607 17163
rect 27685 17085 27690 17163
rect 27602 17080 27690 17085
rect 29936 17160 30256 17216
rect 25936 16896 26256 16920
rect 28360 16916 28600 16940
rect 22810 16711 22946 16716
rect 18810 16632 18946 16637
rect 22810 16637 22815 16711
rect 22941 16637 22946 16711
rect 24360 16700 24600 16724
rect 28360 16724 28384 16916
rect 28576 16724 28600 16916
rect 29936 16920 29960 17160
rect 30224 16920 30256 17160
rect 31602 17163 31690 17168
rect 31602 17085 31607 17163
rect 31685 17085 31690 17163
rect 31602 17080 31690 17085
rect 33936 17160 34256 17216
rect 29936 16896 30256 16920
rect 32360 16916 32600 16940
rect 26810 16711 26946 16716
rect 22810 16632 22946 16637
rect 26810 16637 26815 16711
rect 26941 16637 26946 16711
rect 28360 16700 28600 16724
rect 32360 16724 32384 16916
rect 32576 16724 32600 16916
rect 33936 16920 33960 17160
rect 34224 16920 34256 17160
rect 35602 17163 35690 17168
rect 35602 17085 35607 17163
rect 35685 17085 35690 17163
rect 35602 17080 35690 17085
rect 37936 17160 38256 17216
rect 33936 16896 34256 16920
rect 36360 16916 36600 16940
rect 30810 16711 30946 16716
rect 26810 16632 26946 16637
rect 30810 16637 30815 16711
rect 30941 16637 30946 16711
rect 32360 16700 32600 16724
rect 36360 16724 36384 16916
rect 36576 16724 36600 16916
rect 37936 16920 37960 17160
rect 38224 16920 38256 17160
rect 39602 17163 39690 17168
rect 39602 17085 39607 17163
rect 39685 17085 39690 17163
rect 39602 17080 39690 17085
rect 37936 16896 38256 16920
rect 34810 16711 34946 16716
rect 30810 16632 30946 16637
rect 34810 16637 34815 16711
rect 34941 16637 34946 16711
rect 36360 16700 36600 16724
rect 38810 16711 38946 16716
rect 34810 16632 34946 16637
rect 38810 16637 38815 16711
rect 38941 16637 38946 16711
rect 38810 16632 38946 16637
rect 2338 16573 2518 16574
rect 2338 16395 2339 16573
rect 2517 16395 2518 16573
rect 2338 16394 2518 16395
rect 6338 16573 6518 16574
rect 6338 16395 6339 16573
rect 6517 16395 6518 16573
rect 6338 16394 6518 16395
rect 10338 16573 10518 16574
rect 10338 16395 10339 16573
rect 10517 16395 10518 16573
rect 10338 16394 10518 16395
rect 14338 16573 14518 16574
rect 14338 16395 14339 16573
rect 14517 16395 14518 16573
rect 14338 16394 14518 16395
rect 18338 16573 18518 16574
rect 18338 16395 18339 16573
rect 18517 16395 18518 16573
rect 18338 16394 18518 16395
rect 22338 16573 22518 16574
rect 22338 16395 22339 16573
rect 22517 16395 22518 16573
rect 22338 16394 22518 16395
rect 26338 16573 26518 16574
rect 26338 16395 26339 16573
rect 26517 16395 26518 16573
rect 26338 16394 26518 16395
rect 30338 16573 30518 16574
rect 30338 16395 30339 16573
rect 30517 16395 30518 16573
rect 30338 16394 30518 16395
rect 34338 16573 34518 16574
rect 34338 16395 34339 16573
rect 34517 16395 34518 16573
rect 34338 16394 34518 16395
rect 38338 16573 38518 16574
rect 38338 16395 38339 16573
rect 38517 16395 38518 16573
rect 38338 16394 38518 16395
rect 400 15999 580 16000
rect 400 15821 401 15999
rect 579 15821 580 15999
rect 3734 15996 3740 16002
rect 3780 15996 3786 16002
rect 4400 15999 4580 16000
rect 3728 15990 3734 15996
rect 3786 15990 3792 15996
rect 3728 15944 3734 15950
rect 3786 15944 3792 15950
rect 3734 15938 3740 15944
rect 3780 15938 3786 15944
rect 400 15820 580 15821
rect 4400 15821 4401 15999
rect 4579 15821 4580 15999
rect 7734 15996 7740 16002
rect 7780 15996 7786 16002
rect 8400 15999 8580 16000
rect 7728 15990 7734 15996
rect 7786 15990 7792 15996
rect 7728 15944 7734 15950
rect 7786 15944 7792 15950
rect 7734 15938 7740 15944
rect 7780 15938 7786 15944
rect 4400 15820 4580 15821
rect 8400 15821 8401 15999
rect 8579 15821 8580 15999
rect 11734 15996 11740 16002
rect 11780 15996 11786 16002
rect 12400 15999 12580 16000
rect 11728 15990 11734 15996
rect 11786 15990 11792 15996
rect 11728 15944 11734 15950
rect 11786 15944 11792 15950
rect 11734 15938 11740 15944
rect 11780 15938 11786 15944
rect 8400 15820 8580 15821
rect 12400 15821 12401 15999
rect 12579 15821 12580 15999
rect 15734 15996 15740 16002
rect 15780 15996 15786 16002
rect 16400 15999 16580 16000
rect 15728 15990 15734 15996
rect 15786 15990 15792 15996
rect 15728 15944 15734 15950
rect 15786 15944 15792 15950
rect 15734 15938 15740 15944
rect 15780 15938 15786 15944
rect 12400 15820 12580 15821
rect 16400 15821 16401 15999
rect 16579 15821 16580 15999
rect 19734 15996 19740 16002
rect 19780 15996 19786 16002
rect 20400 15999 20580 16000
rect 19728 15990 19734 15996
rect 19786 15990 19792 15996
rect 19728 15944 19734 15950
rect 19786 15944 19792 15950
rect 19734 15938 19740 15944
rect 19780 15938 19786 15944
rect 16400 15820 16580 15821
rect 20400 15821 20401 15999
rect 20579 15821 20580 15999
rect 23734 15996 23740 16002
rect 23780 15996 23786 16002
rect 24400 15999 24580 16000
rect 23728 15990 23734 15996
rect 23786 15990 23792 15996
rect 23728 15944 23734 15950
rect 23786 15944 23792 15950
rect 23734 15938 23740 15944
rect 23780 15938 23786 15944
rect 20400 15820 20580 15821
rect 24400 15821 24401 15999
rect 24579 15821 24580 15999
rect 27734 15996 27740 16002
rect 27780 15996 27786 16002
rect 28400 15999 28580 16000
rect 27728 15990 27734 15996
rect 27786 15990 27792 15996
rect 27728 15944 27734 15950
rect 27786 15944 27792 15950
rect 27734 15938 27740 15944
rect 27780 15938 27786 15944
rect 24400 15820 24580 15821
rect 28400 15821 28401 15999
rect 28579 15821 28580 15999
rect 31734 15996 31740 16002
rect 31780 15996 31786 16002
rect 32400 15999 32580 16000
rect 31728 15990 31734 15996
rect 31786 15990 31792 15996
rect 31728 15944 31734 15950
rect 31786 15944 31792 15950
rect 31734 15938 31740 15944
rect 31780 15938 31786 15944
rect 28400 15820 28580 15821
rect 32400 15821 32401 15999
rect 32579 15821 32580 15999
rect 35734 15996 35740 16002
rect 35780 15996 35786 16002
rect 36400 15999 36580 16000
rect 35728 15990 35734 15996
rect 35786 15990 35792 15996
rect 35728 15944 35734 15950
rect 35786 15944 35792 15950
rect 35734 15938 35740 15944
rect 35780 15938 35786 15944
rect 32400 15820 32580 15821
rect 36400 15821 36401 15999
rect 36579 15821 36580 15999
rect 39734 15996 39740 16002
rect 39780 15996 39786 16002
rect 39728 15990 39734 15996
rect 39786 15990 39792 15996
rect 39728 15944 39734 15950
rect 39786 15944 39792 15950
rect 39734 15938 39740 15944
rect 39780 15938 39786 15944
rect 36400 15820 36580 15821
rect 3262 15808 3268 15814
rect 3308 15808 3314 15814
rect 7262 15808 7268 15814
rect 7308 15808 7314 15814
rect 11262 15808 11268 15814
rect 11308 15808 11314 15814
rect 15262 15808 15268 15814
rect 15308 15808 15314 15814
rect 19262 15808 19268 15814
rect 19308 15808 19314 15814
rect 23262 15808 23268 15814
rect 23308 15808 23314 15814
rect 27262 15808 27268 15814
rect 27308 15808 27314 15814
rect 31262 15808 31268 15814
rect 31308 15808 31314 15814
rect 35262 15808 35268 15814
rect 35308 15808 35314 15814
rect 39262 15808 39268 15814
rect 39308 15808 39314 15814
rect 3256 15802 3262 15808
rect 3314 15802 3320 15808
rect 7256 15802 7262 15808
rect 7314 15802 7320 15808
rect 11256 15802 11262 15808
rect 11314 15802 11320 15808
rect 15256 15802 15262 15808
rect 15314 15802 15320 15808
rect 19256 15802 19262 15808
rect 19314 15802 19320 15808
rect 23256 15802 23262 15808
rect 23314 15802 23320 15808
rect 27256 15802 27262 15808
rect 27314 15802 27320 15808
rect 31256 15802 31262 15808
rect 31314 15802 31320 15808
rect 35256 15802 35262 15808
rect 35314 15802 35320 15808
rect 39256 15802 39262 15808
rect 39314 15802 39320 15808
rect 3256 15756 3262 15762
rect 3314 15756 3320 15762
rect 7256 15756 7262 15762
rect 7314 15756 7320 15762
rect 11256 15756 11262 15762
rect 11314 15756 11320 15762
rect 15256 15756 15262 15762
rect 15314 15756 15320 15762
rect 19256 15756 19262 15762
rect 19314 15756 19320 15762
rect 23256 15756 23262 15762
rect 23314 15756 23320 15762
rect 27256 15756 27262 15762
rect 27314 15756 27320 15762
rect 31256 15756 31262 15762
rect 31314 15756 31320 15762
rect 35256 15756 35262 15762
rect 35314 15756 35320 15762
rect 39256 15756 39262 15762
rect 39314 15756 39320 15762
rect 3262 15750 3268 15756
rect 3308 15750 3314 15756
rect 7262 15750 7268 15756
rect 7308 15750 7314 15756
rect 11262 15750 11268 15756
rect 11308 15750 11314 15756
rect 15262 15750 15268 15756
rect 15308 15750 15314 15756
rect 19262 15750 19268 15756
rect 19308 15750 19314 15756
rect 23262 15750 23268 15756
rect 23308 15750 23314 15756
rect 27262 15750 27268 15756
rect 27308 15750 27314 15756
rect 31262 15750 31268 15756
rect 31308 15750 31314 15756
rect 35262 15750 35268 15756
rect 35308 15750 35314 15756
rect 39262 15750 39268 15756
rect 39308 15750 39314 15756
rect 2240 15296 2480 15320
rect 2240 15104 2264 15296
rect 2456 15104 2480 15296
rect 2240 15080 2480 15104
rect 6240 15296 6480 15320
rect 6240 15104 6264 15296
rect 6456 15104 6480 15296
rect 6240 15080 6480 15104
rect 10240 15296 10480 15320
rect 10240 15104 10264 15296
rect 10456 15104 10480 15296
rect 10240 15080 10480 15104
rect 14240 15296 14480 15320
rect 14240 15104 14264 15296
rect 14456 15104 14480 15296
rect 14240 15080 14480 15104
rect 18240 15296 18480 15320
rect 18240 15104 18264 15296
rect 18456 15104 18480 15296
rect 18240 15080 18480 15104
rect 22240 15296 22480 15320
rect 22240 15104 22264 15296
rect 22456 15104 22480 15296
rect 22240 15080 22480 15104
rect 26240 15296 26480 15320
rect 26240 15104 26264 15296
rect 26456 15104 26480 15296
rect 26240 15080 26480 15104
rect 30240 15296 30480 15320
rect 30240 15104 30264 15296
rect 30456 15104 30480 15296
rect 30240 15080 30480 15104
rect 34240 15296 34480 15320
rect 34240 15104 34264 15296
rect 34456 15104 34480 15296
rect 34240 15080 34480 15104
rect 38240 15296 38480 15320
rect 38240 15104 38264 15296
rect 38456 15104 38480 15296
rect 38240 15080 38480 15104
rect 2240 14596 2480 14620
rect 2240 14536 2264 14596
rect 2456 14536 2480 14596
rect 2240 14380 2480 14536
rect 6240 14596 6480 14620
rect 6240 14536 6264 14596
rect 6456 14536 6480 14596
rect 6240 14380 6480 14536
rect 10240 14596 10480 14620
rect 10240 14536 10264 14596
rect 10456 14536 10480 14596
rect 10240 14380 10480 14536
rect 14240 14596 14480 14620
rect 14240 14536 14264 14596
rect 14456 14536 14480 14596
rect 14240 14380 14480 14536
rect 18240 14596 18480 14620
rect 18240 14536 18264 14596
rect 18456 14536 18480 14596
rect 18240 14380 18480 14536
rect 22240 14596 22480 14620
rect 22240 14536 22264 14596
rect 22456 14536 22480 14596
rect 22240 14380 22480 14536
rect 26240 14596 26480 14620
rect 26240 14536 26264 14596
rect 26456 14536 26480 14596
rect 26240 14380 26480 14536
rect 30240 14596 30480 14620
rect 30240 14536 30264 14596
rect 30456 14536 30480 14596
rect 30240 14380 30480 14536
rect 34240 14596 34480 14620
rect 34240 14536 34264 14596
rect 34456 14536 34480 14596
rect 34240 14380 34480 14536
rect 38240 14596 38480 14620
rect 38240 14536 38264 14596
rect 38456 14536 38480 14596
rect 38240 14380 38480 14536
rect 1936 14160 2256 14216
rect 360 13916 600 13940
rect 360 13724 384 13916
rect 576 13724 600 13916
rect 1936 13920 1960 14160
rect 2224 13920 2256 14160
rect 3602 14163 3690 14168
rect 3602 14085 3607 14163
rect 3685 14085 3690 14163
rect 3602 14080 3690 14085
rect 5936 14160 6256 14216
rect 1936 13896 2256 13920
rect 4360 13916 4600 13940
rect 360 13700 600 13724
rect 4360 13724 4384 13916
rect 4576 13724 4600 13916
rect 5936 13920 5960 14160
rect 6224 13920 6256 14160
rect 7602 14163 7690 14168
rect 7602 14085 7607 14163
rect 7685 14085 7690 14163
rect 7602 14080 7690 14085
rect 9936 14160 10256 14216
rect 5936 13896 6256 13920
rect 8360 13916 8600 13940
rect 2810 13711 2946 13716
rect 2810 13637 2815 13711
rect 2941 13637 2946 13711
rect 4360 13700 4600 13724
rect 8360 13724 8384 13916
rect 8576 13724 8600 13916
rect 9936 13920 9960 14160
rect 10224 13920 10256 14160
rect 11602 14163 11690 14168
rect 11602 14085 11607 14163
rect 11685 14085 11690 14163
rect 11602 14080 11690 14085
rect 13936 14160 14256 14216
rect 9936 13896 10256 13920
rect 12360 13916 12600 13940
rect 6810 13711 6946 13716
rect 2810 13632 2946 13637
rect 6810 13637 6815 13711
rect 6941 13637 6946 13711
rect 8360 13700 8600 13724
rect 12360 13724 12384 13916
rect 12576 13724 12600 13916
rect 13936 13920 13960 14160
rect 14224 13920 14256 14160
rect 15602 14163 15690 14168
rect 15602 14085 15607 14163
rect 15685 14085 15690 14163
rect 15602 14080 15690 14085
rect 17936 14160 18256 14216
rect 13936 13896 14256 13920
rect 16360 13916 16600 13940
rect 10810 13711 10946 13716
rect 6810 13632 6946 13637
rect 10810 13637 10815 13711
rect 10941 13637 10946 13711
rect 12360 13700 12600 13724
rect 16360 13724 16384 13916
rect 16576 13724 16600 13916
rect 17936 13920 17960 14160
rect 18224 13920 18256 14160
rect 19602 14163 19690 14168
rect 19602 14085 19607 14163
rect 19685 14085 19690 14163
rect 19602 14080 19690 14085
rect 21936 14160 22256 14216
rect 17936 13896 18256 13920
rect 20360 13916 20600 13940
rect 14810 13711 14946 13716
rect 10810 13632 10946 13637
rect 14810 13637 14815 13711
rect 14941 13637 14946 13711
rect 16360 13700 16600 13724
rect 20360 13724 20384 13916
rect 20576 13724 20600 13916
rect 21936 13920 21960 14160
rect 22224 13920 22256 14160
rect 23602 14163 23690 14168
rect 23602 14085 23607 14163
rect 23685 14085 23690 14163
rect 23602 14080 23690 14085
rect 25936 14160 26256 14216
rect 21936 13896 22256 13920
rect 24360 13916 24600 13940
rect 18810 13711 18946 13716
rect 14810 13632 14946 13637
rect 18810 13637 18815 13711
rect 18941 13637 18946 13711
rect 20360 13700 20600 13724
rect 24360 13724 24384 13916
rect 24576 13724 24600 13916
rect 25936 13920 25960 14160
rect 26224 13920 26256 14160
rect 27602 14163 27690 14168
rect 27602 14085 27607 14163
rect 27685 14085 27690 14163
rect 27602 14080 27690 14085
rect 29936 14160 30256 14216
rect 25936 13896 26256 13920
rect 28360 13916 28600 13940
rect 22810 13711 22946 13716
rect 18810 13632 18946 13637
rect 22810 13637 22815 13711
rect 22941 13637 22946 13711
rect 24360 13700 24600 13724
rect 28360 13724 28384 13916
rect 28576 13724 28600 13916
rect 29936 13920 29960 14160
rect 30224 13920 30256 14160
rect 31602 14163 31690 14168
rect 31602 14085 31607 14163
rect 31685 14085 31690 14163
rect 31602 14080 31690 14085
rect 33936 14160 34256 14216
rect 29936 13896 30256 13920
rect 32360 13916 32600 13940
rect 26810 13711 26946 13716
rect 22810 13632 22946 13637
rect 26810 13637 26815 13711
rect 26941 13637 26946 13711
rect 28360 13700 28600 13724
rect 32360 13724 32384 13916
rect 32576 13724 32600 13916
rect 33936 13920 33960 14160
rect 34224 13920 34256 14160
rect 35602 14163 35690 14168
rect 35602 14085 35607 14163
rect 35685 14085 35690 14163
rect 35602 14080 35690 14085
rect 37936 14160 38256 14216
rect 33936 13896 34256 13920
rect 36360 13916 36600 13940
rect 30810 13711 30946 13716
rect 26810 13632 26946 13637
rect 30810 13637 30815 13711
rect 30941 13637 30946 13711
rect 32360 13700 32600 13724
rect 36360 13724 36384 13916
rect 36576 13724 36600 13916
rect 37936 13920 37960 14160
rect 38224 13920 38256 14160
rect 39602 14163 39690 14168
rect 39602 14085 39607 14163
rect 39685 14085 39690 14163
rect 39602 14080 39690 14085
rect 37936 13896 38256 13920
rect 34810 13711 34946 13716
rect 30810 13632 30946 13637
rect 34810 13637 34815 13711
rect 34941 13637 34946 13711
rect 36360 13700 36600 13724
rect 38810 13711 38946 13716
rect 34810 13632 34946 13637
rect 38810 13637 38815 13711
rect 38941 13637 38946 13711
rect 38810 13632 38946 13637
rect 2338 13573 2518 13574
rect 2338 13395 2339 13573
rect 2517 13395 2518 13573
rect 2338 13394 2518 13395
rect 6338 13573 6518 13574
rect 6338 13395 6339 13573
rect 6517 13395 6518 13573
rect 6338 13394 6518 13395
rect 10338 13573 10518 13574
rect 10338 13395 10339 13573
rect 10517 13395 10518 13573
rect 10338 13394 10518 13395
rect 14338 13573 14518 13574
rect 14338 13395 14339 13573
rect 14517 13395 14518 13573
rect 14338 13394 14518 13395
rect 18338 13573 18518 13574
rect 18338 13395 18339 13573
rect 18517 13395 18518 13573
rect 18338 13394 18518 13395
rect 22338 13573 22518 13574
rect 22338 13395 22339 13573
rect 22517 13395 22518 13573
rect 22338 13394 22518 13395
rect 26338 13573 26518 13574
rect 26338 13395 26339 13573
rect 26517 13395 26518 13573
rect 26338 13394 26518 13395
rect 30338 13573 30518 13574
rect 30338 13395 30339 13573
rect 30517 13395 30518 13573
rect 30338 13394 30518 13395
rect 34338 13573 34518 13574
rect 34338 13395 34339 13573
rect 34517 13395 34518 13573
rect 34338 13394 34518 13395
rect 38338 13573 38518 13574
rect 38338 13395 38339 13573
rect 38517 13395 38518 13573
rect 38338 13394 38518 13395
rect 400 12999 580 13000
rect 400 12821 401 12999
rect 579 12821 580 12999
rect 3734 12996 3740 13002
rect 3780 12996 3786 13002
rect 4400 12999 4580 13000
rect 3728 12990 3734 12996
rect 3786 12990 3792 12996
rect 3728 12944 3734 12950
rect 3786 12944 3792 12950
rect 3734 12938 3740 12944
rect 3780 12938 3786 12944
rect 400 12820 580 12821
rect 4400 12821 4401 12999
rect 4579 12821 4580 12999
rect 7734 12996 7740 13002
rect 7780 12996 7786 13002
rect 8400 12999 8580 13000
rect 7728 12990 7734 12996
rect 7786 12990 7792 12996
rect 7728 12944 7734 12950
rect 7786 12944 7792 12950
rect 7734 12938 7740 12944
rect 7780 12938 7786 12944
rect 4400 12820 4580 12821
rect 8400 12821 8401 12999
rect 8579 12821 8580 12999
rect 11734 12996 11740 13002
rect 11780 12996 11786 13002
rect 12400 12999 12580 13000
rect 11728 12990 11734 12996
rect 11786 12990 11792 12996
rect 11728 12944 11734 12950
rect 11786 12944 11792 12950
rect 11734 12938 11740 12944
rect 11780 12938 11786 12944
rect 8400 12820 8580 12821
rect 12400 12821 12401 12999
rect 12579 12821 12580 12999
rect 15734 12996 15740 13002
rect 15780 12996 15786 13002
rect 16400 12999 16580 13000
rect 15728 12990 15734 12996
rect 15786 12990 15792 12996
rect 15728 12944 15734 12950
rect 15786 12944 15792 12950
rect 15734 12938 15740 12944
rect 15780 12938 15786 12944
rect 12400 12820 12580 12821
rect 16400 12821 16401 12999
rect 16579 12821 16580 12999
rect 19734 12996 19740 13002
rect 19780 12996 19786 13002
rect 20400 12999 20580 13000
rect 19728 12990 19734 12996
rect 19786 12990 19792 12996
rect 19728 12944 19734 12950
rect 19786 12944 19792 12950
rect 19734 12938 19740 12944
rect 19780 12938 19786 12944
rect 16400 12820 16580 12821
rect 20400 12821 20401 12999
rect 20579 12821 20580 12999
rect 23734 12996 23740 13002
rect 23780 12996 23786 13002
rect 24400 12999 24580 13000
rect 23728 12990 23734 12996
rect 23786 12990 23792 12996
rect 23728 12944 23734 12950
rect 23786 12944 23792 12950
rect 23734 12938 23740 12944
rect 23780 12938 23786 12944
rect 20400 12820 20580 12821
rect 24400 12821 24401 12999
rect 24579 12821 24580 12999
rect 27734 12996 27740 13002
rect 27780 12996 27786 13002
rect 28400 12999 28580 13000
rect 27728 12990 27734 12996
rect 27786 12990 27792 12996
rect 27728 12944 27734 12950
rect 27786 12944 27792 12950
rect 27734 12938 27740 12944
rect 27780 12938 27786 12944
rect 24400 12820 24580 12821
rect 28400 12821 28401 12999
rect 28579 12821 28580 12999
rect 31734 12996 31740 13002
rect 31780 12996 31786 13002
rect 32400 12999 32580 13000
rect 31728 12990 31734 12996
rect 31786 12990 31792 12996
rect 31728 12944 31734 12950
rect 31786 12944 31792 12950
rect 31734 12938 31740 12944
rect 31780 12938 31786 12944
rect 28400 12820 28580 12821
rect 32400 12821 32401 12999
rect 32579 12821 32580 12999
rect 35734 12996 35740 13002
rect 35780 12996 35786 13002
rect 36400 12999 36580 13000
rect 35728 12990 35734 12996
rect 35786 12990 35792 12996
rect 35728 12944 35734 12950
rect 35786 12944 35792 12950
rect 35734 12938 35740 12944
rect 35780 12938 35786 12944
rect 32400 12820 32580 12821
rect 36400 12821 36401 12999
rect 36579 12821 36580 12999
rect 39734 12996 39740 13002
rect 39780 12996 39786 13002
rect 39728 12990 39734 12996
rect 39786 12990 39792 12996
rect 39728 12944 39734 12950
rect 39786 12944 39792 12950
rect 39734 12938 39740 12944
rect 39780 12938 39786 12944
rect 36400 12820 36580 12821
rect 3262 12808 3268 12814
rect 3308 12808 3314 12814
rect 7262 12808 7268 12814
rect 7308 12808 7314 12814
rect 11262 12808 11268 12814
rect 11308 12808 11314 12814
rect 15262 12808 15268 12814
rect 15308 12808 15314 12814
rect 19262 12808 19268 12814
rect 19308 12808 19314 12814
rect 23262 12808 23268 12814
rect 23308 12808 23314 12814
rect 27262 12808 27268 12814
rect 27308 12808 27314 12814
rect 31262 12808 31268 12814
rect 31308 12808 31314 12814
rect 35262 12808 35268 12814
rect 35308 12808 35314 12814
rect 39262 12808 39268 12814
rect 39308 12808 39314 12814
rect 3256 12802 3262 12808
rect 3314 12802 3320 12808
rect 7256 12802 7262 12808
rect 7314 12802 7320 12808
rect 11256 12802 11262 12808
rect 11314 12802 11320 12808
rect 15256 12802 15262 12808
rect 15314 12802 15320 12808
rect 19256 12802 19262 12808
rect 19314 12802 19320 12808
rect 23256 12802 23262 12808
rect 23314 12802 23320 12808
rect 27256 12802 27262 12808
rect 27314 12802 27320 12808
rect 31256 12802 31262 12808
rect 31314 12802 31320 12808
rect 35256 12802 35262 12808
rect 35314 12802 35320 12808
rect 39256 12802 39262 12808
rect 39314 12802 39320 12808
rect 3256 12756 3262 12762
rect 3314 12756 3320 12762
rect 7256 12756 7262 12762
rect 7314 12756 7320 12762
rect 11256 12756 11262 12762
rect 11314 12756 11320 12762
rect 15256 12756 15262 12762
rect 15314 12756 15320 12762
rect 19256 12756 19262 12762
rect 19314 12756 19320 12762
rect 23256 12756 23262 12762
rect 23314 12756 23320 12762
rect 27256 12756 27262 12762
rect 27314 12756 27320 12762
rect 31256 12756 31262 12762
rect 31314 12756 31320 12762
rect 35256 12756 35262 12762
rect 35314 12756 35320 12762
rect 39256 12756 39262 12762
rect 39314 12756 39320 12762
rect 3262 12750 3268 12756
rect 3308 12750 3314 12756
rect 7262 12750 7268 12756
rect 7308 12750 7314 12756
rect 11262 12750 11268 12756
rect 11308 12750 11314 12756
rect 15262 12750 15268 12756
rect 15308 12750 15314 12756
rect 19262 12750 19268 12756
rect 19308 12750 19314 12756
rect 23262 12750 23268 12756
rect 23308 12750 23314 12756
rect 27262 12750 27268 12756
rect 27308 12750 27314 12756
rect 31262 12750 31268 12756
rect 31308 12750 31314 12756
rect 35262 12750 35268 12756
rect 35308 12750 35314 12756
rect 39262 12750 39268 12756
rect 39308 12750 39314 12756
rect 2240 12296 2480 12320
rect 2240 12104 2264 12296
rect 2456 12104 2480 12296
rect 2240 12080 2480 12104
rect 6240 12296 6480 12320
rect 6240 12104 6264 12296
rect 6456 12104 6480 12296
rect 6240 12080 6480 12104
rect 10240 12296 10480 12320
rect 10240 12104 10264 12296
rect 10456 12104 10480 12296
rect 10240 12080 10480 12104
rect 14240 12296 14480 12320
rect 14240 12104 14264 12296
rect 14456 12104 14480 12296
rect 14240 12080 14480 12104
rect 18240 12296 18480 12320
rect 18240 12104 18264 12296
rect 18456 12104 18480 12296
rect 18240 12080 18480 12104
rect 22240 12296 22480 12320
rect 22240 12104 22264 12296
rect 22456 12104 22480 12296
rect 22240 12080 22480 12104
rect 26240 12296 26480 12320
rect 26240 12104 26264 12296
rect 26456 12104 26480 12296
rect 26240 12080 26480 12104
rect 30240 12296 30480 12320
rect 30240 12104 30264 12296
rect 30456 12104 30480 12296
rect 30240 12080 30480 12104
rect 34240 12296 34480 12320
rect 34240 12104 34264 12296
rect 34456 12104 34480 12296
rect 34240 12080 34480 12104
rect 38240 12296 38480 12320
rect 38240 12104 38264 12296
rect 38456 12104 38480 12296
rect 38240 12080 38480 12104
rect 2240 11596 2480 11620
rect 2240 11536 2264 11596
rect 2456 11536 2480 11596
rect 2240 11380 2480 11536
rect 6240 11596 6480 11620
rect 6240 11536 6264 11596
rect 6456 11536 6480 11596
rect 6240 11380 6480 11536
rect 10240 11596 10480 11620
rect 10240 11536 10264 11596
rect 10456 11536 10480 11596
rect 10240 11380 10480 11536
rect 14240 11596 14480 11620
rect 14240 11536 14264 11596
rect 14456 11536 14480 11596
rect 14240 11380 14480 11536
rect 18240 11596 18480 11620
rect 18240 11536 18264 11596
rect 18456 11536 18480 11596
rect 18240 11380 18480 11536
rect 22240 11596 22480 11620
rect 22240 11536 22264 11596
rect 22456 11536 22480 11596
rect 22240 11380 22480 11536
rect 26240 11596 26480 11620
rect 26240 11536 26264 11596
rect 26456 11536 26480 11596
rect 26240 11380 26480 11536
rect 30240 11596 30480 11620
rect 30240 11536 30264 11596
rect 30456 11536 30480 11596
rect 30240 11380 30480 11536
rect 34240 11596 34480 11620
rect 34240 11536 34264 11596
rect 34456 11536 34480 11596
rect 34240 11380 34480 11536
rect 38240 11596 38480 11620
rect 38240 11536 38264 11596
rect 38456 11536 38480 11596
rect 38240 11380 38480 11536
rect 1936 11160 2256 11216
rect 360 10916 600 10940
rect 360 10724 384 10916
rect 576 10724 600 10916
rect 1936 10920 1960 11160
rect 2224 10920 2256 11160
rect 3602 11163 3690 11168
rect 3602 11085 3607 11163
rect 3685 11085 3690 11163
rect 3602 11080 3690 11085
rect 5936 11160 6256 11216
rect 1936 10896 2256 10920
rect 4360 10916 4600 10940
rect 360 10700 600 10724
rect 4360 10724 4384 10916
rect 4576 10724 4600 10916
rect 5936 10920 5960 11160
rect 6224 10920 6256 11160
rect 7602 11163 7690 11168
rect 7602 11085 7607 11163
rect 7685 11085 7690 11163
rect 7602 11080 7690 11085
rect 9936 11160 10256 11216
rect 5936 10896 6256 10920
rect 8360 10916 8600 10940
rect 2810 10711 2946 10716
rect 2810 10637 2815 10711
rect 2941 10637 2946 10711
rect 4360 10700 4600 10724
rect 8360 10724 8384 10916
rect 8576 10724 8600 10916
rect 9936 10920 9960 11160
rect 10224 10920 10256 11160
rect 11602 11163 11690 11168
rect 11602 11085 11607 11163
rect 11685 11085 11690 11163
rect 11602 11080 11690 11085
rect 13936 11160 14256 11216
rect 9936 10896 10256 10920
rect 12360 10916 12600 10940
rect 6810 10711 6946 10716
rect 2810 10632 2946 10637
rect 6810 10637 6815 10711
rect 6941 10637 6946 10711
rect 8360 10700 8600 10724
rect 12360 10724 12384 10916
rect 12576 10724 12600 10916
rect 13936 10920 13960 11160
rect 14224 10920 14256 11160
rect 15602 11163 15690 11168
rect 15602 11085 15607 11163
rect 15685 11085 15690 11163
rect 15602 11080 15690 11085
rect 17936 11160 18256 11216
rect 13936 10896 14256 10920
rect 16360 10916 16600 10940
rect 10810 10711 10946 10716
rect 6810 10632 6946 10637
rect 10810 10637 10815 10711
rect 10941 10637 10946 10711
rect 12360 10700 12600 10724
rect 16360 10724 16384 10916
rect 16576 10724 16600 10916
rect 17936 10920 17960 11160
rect 18224 10920 18256 11160
rect 19602 11163 19690 11168
rect 19602 11085 19607 11163
rect 19685 11085 19690 11163
rect 19602 11080 19690 11085
rect 21936 11160 22256 11216
rect 17936 10896 18256 10920
rect 20360 10916 20600 10940
rect 14810 10711 14946 10716
rect 10810 10632 10946 10637
rect 14810 10637 14815 10711
rect 14941 10637 14946 10711
rect 16360 10700 16600 10724
rect 20360 10724 20384 10916
rect 20576 10724 20600 10916
rect 21936 10920 21960 11160
rect 22224 10920 22256 11160
rect 23602 11163 23690 11168
rect 23602 11085 23607 11163
rect 23685 11085 23690 11163
rect 23602 11080 23690 11085
rect 25936 11160 26256 11216
rect 21936 10896 22256 10920
rect 24360 10916 24600 10940
rect 18810 10711 18946 10716
rect 14810 10632 14946 10637
rect 18810 10637 18815 10711
rect 18941 10637 18946 10711
rect 20360 10700 20600 10724
rect 24360 10724 24384 10916
rect 24576 10724 24600 10916
rect 25936 10920 25960 11160
rect 26224 10920 26256 11160
rect 27602 11163 27690 11168
rect 27602 11085 27607 11163
rect 27685 11085 27690 11163
rect 27602 11080 27690 11085
rect 29936 11160 30256 11216
rect 25936 10896 26256 10920
rect 28360 10916 28600 10940
rect 22810 10711 22946 10716
rect 18810 10632 18946 10637
rect 22810 10637 22815 10711
rect 22941 10637 22946 10711
rect 24360 10700 24600 10724
rect 28360 10724 28384 10916
rect 28576 10724 28600 10916
rect 29936 10920 29960 11160
rect 30224 10920 30256 11160
rect 31602 11163 31690 11168
rect 31602 11085 31607 11163
rect 31685 11085 31690 11163
rect 31602 11080 31690 11085
rect 33936 11160 34256 11216
rect 29936 10896 30256 10920
rect 32360 10916 32600 10940
rect 26810 10711 26946 10716
rect 22810 10632 22946 10637
rect 26810 10637 26815 10711
rect 26941 10637 26946 10711
rect 28360 10700 28600 10724
rect 32360 10724 32384 10916
rect 32576 10724 32600 10916
rect 33936 10920 33960 11160
rect 34224 10920 34256 11160
rect 35602 11163 35690 11168
rect 35602 11085 35607 11163
rect 35685 11085 35690 11163
rect 35602 11080 35690 11085
rect 37936 11160 38256 11216
rect 33936 10896 34256 10920
rect 36360 10916 36600 10940
rect 30810 10711 30946 10716
rect 26810 10632 26946 10637
rect 30810 10637 30815 10711
rect 30941 10637 30946 10711
rect 32360 10700 32600 10724
rect 36360 10724 36384 10916
rect 36576 10724 36600 10916
rect 37936 10920 37960 11160
rect 38224 10920 38256 11160
rect 39602 11163 39690 11168
rect 39602 11085 39607 11163
rect 39685 11085 39690 11163
rect 39602 11080 39690 11085
rect 37936 10896 38256 10920
rect 34810 10711 34946 10716
rect 30810 10632 30946 10637
rect 34810 10637 34815 10711
rect 34941 10637 34946 10711
rect 36360 10700 36600 10724
rect 38810 10711 38946 10716
rect 34810 10632 34946 10637
rect 38810 10637 38815 10711
rect 38941 10637 38946 10711
rect 38810 10632 38946 10637
rect 2338 10573 2518 10574
rect 2338 10395 2339 10573
rect 2517 10395 2518 10573
rect 2338 10394 2518 10395
rect 6338 10573 6518 10574
rect 6338 10395 6339 10573
rect 6517 10395 6518 10573
rect 6338 10394 6518 10395
rect 10338 10573 10518 10574
rect 10338 10395 10339 10573
rect 10517 10395 10518 10573
rect 10338 10394 10518 10395
rect 14338 10573 14518 10574
rect 14338 10395 14339 10573
rect 14517 10395 14518 10573
rect 14338 10394 14518 10395
rect 18338 10573 18518 10574
rect 18338 10395 18339 10573
rect 18517 10395 18518 10573
rect 18338 10394 18518 10395
rect 22338 10573 22518 10574
rect 22338 10395 22339 10573
rect 22517 10395 22518 10573
rect 22338 10394 22518 10395
rect 26338 10573 26518 10574
rect 26338 10395 26339 10573
rect 26517 10395 26518 10573
rect 26338 10394 26518 10395
rect 30338 10573 30518 10574
rect 30338 10395 30339 10573
rect 30517 10395 30518 10573
rect 30338 10394 30518 10395
rect 34338 10573 34518 10574
rect 34338 10395 34339 10573
rect 34517 10395 34518 10573
rect 34338 10394 34518 10395
rect 38338 10573 38518 10574
rect 38338 10395 38339 10573
rect 38517 10395 38518 10573
rect 38338 10394 38518 10395
rect 400 9999 580 10000
rect 400 9821 401 9999
rect 579 9821 580 9999
rect 3734 9996 3740 10002
rect 3780 9996 3786 10002
rect 4400 9999 4580 10000
rect 3728 9990 3734 9996
rect 3786 9990 3792 9996
rect 3728 9944 3734 9950
rect 3786 9944 3792 9950
rect 3734 9938 3740 9944
rect 3780 9938 3786 9944
rect 400 9820 580 9821
rect 4400 9821 4401 9999
rect 4579 9821 4580 9999
rect 7734 9996 7740 10002
rect 7780 9996 7786 10002
rect 8400 9999 8580 10000
rect 7728 9990 7734 9996
rect 7786 9990 7792 9996
rect 7728 9944 7734 9950
rect 7786 9944 7792 9950
rect 7734 9938 7740 9944
rect 7780 9938 7786 9944
rect 4400 9820 4580 9821
rect 8400 9821 8401 9999
rect 8579 9821 8580 9999
rect 11734 9996 11740 10002
rect 11780 9996 11786 10002
rect 12400 9999 12580 10000
rect 11728 9990 11734 9996
rect 11786 9990 11792 9996
rect 11728 9944 11734 9950
rect 11786 9944 11792 9950
rect 11734 9938 11740 9944
rect 11780 9938 11786 9944
rect 8400 9820 8580 9821
rect 12400 9821 12401 9999
rect 12579 9821 12580 9999
rect 15734 9996 15740 10002
rect 15780 9996 15786 10002
rect 16400 9999 16580 10000
rect 15728 9990 15734 9996
rect 15786 9990 15792 9996
rect 15728 9944 15734 9950
rect 15786 9944 15792 9950
rect 15734 9938 15740 9944
rect 15780 9938 15786 9944
rect 12400 9820 12580 9821
rect 16400 9821 16401 9999
rect 16579 9821 16580 9999
rect 19734 9996 19740 10002
rect 19780 9996 19786 10002
rect 20400 9999 20580 10000
rect 19728 9990 19734 9996
rect 19786 9990 19792 9996
rect 19728 9944 19734 9950
rect 19786 9944 19792 9950
rect 19734 9938 19740 9944
rect 19780 9938 19786 9944
rect 16400 9820 16580 9821
rect 20400 9821 20401 9999
rect 20579 9821 20580 9999
rect 23734 9996 23740 10002
rect 23780 9996 23786 10002
rect 24400 9999 24580 10000
rect 23728 9990 23734 9996
rect 23786 9990 23792 9996
rect 23728 9944 23734 9950
rect 23786 9944 23792 9950
rect 23734 9938 23740 9944
rect 23780 9938 23786 9944
rect 20400 9820 20580 9821
rect 24400 9821 24401 9999
rect 24579 9821 24580 9999
rect 27734 9996 27740 10002
rect 27780 9996 27786 10002
rect 28400 9999 28580 10000
rect 27728 9990 27734 9996
rect 27786 9990 27792 9996
rect 27728 9944 27734 9950
rect 27786 9944 27792 9950
rect 27734 9938 27740 9944
rect 27780 9938 27786 9944
rect 24400 9820 24580 9821
rect 28400 9821 28401 9999
rect 28579 9821 28580 9999
rect 31734 9996 31740 10002
rect 31780 9996 31786 10002
rect 32400 9999 32580 10000
rect 31728 9990 31734 9996
rect 31786 9990 31792 9996
rect 31728 9944 31734 9950
rect 31786 9944 31792 9950
rect 31734 9938 31740 9944
rect 31780 9938 31786 9944
rect 28400 9820 28580 9821
rect 32400 9821 32401 9999
rect 32579 9821 32580 9999
rect 35734 9996 35740 10002
rect 35780 9996 35786 10002
rect 36400 9999 36580 10000
rect 35728 9990 35734 9996
rect 35786 9990 35792 9996
rect 35728 9944 35734 9950
rect 35786 9944 35792 9950
rect 35734 9938 35740 9944
rect 35780 9938 35786 9944
rect 32400 9820 32580 9821
rect 36400 9821 36401 9999
rect 36579 9821 36580 9999
rect 39734 9996 39740 10002
rect 39780 9996 39786 10002
rect 39728 9990 39734 9996
rect 39786 9990 39792 9996
rect 39728 9944 39734 9950
rect 39786 9944 39792 9950
rect 39734 9938 39740 9944
rect 39780 9938 39786 9944
rect 36400 9820 36580 9821
rect 3262 9808 3268 9814
rect 3308 9808 3314 9814
rect 7262 9808 7268 9814
rect 7308 9808 7314 9814
rect 11262 9808 11268 9814
rect 11308 9808 11314 9814
rect 15262 9808 15268 9814
rect 15308 9808 15314 9814
rect 19262 9808 19268 9814
rect 19308 9808 19314 9814
rect 23262 9808 23268 9814
rect 23308 9808 23314 9814
rect 27262 9808 27268 9814
rect 27308 9808 27314 9814
rect 31262 9808 31268 9814
rect 31308 9808 31314 9814
rect 35262 9808 35268 9814
rect 35308 9808 35314 9814
rect 39262 9808 39268 9814
rect 39308 9808 39314 9814
rect 3256 9802 3262 9808
rect 3314 9802 3320 9808
rect 7256 9802 7262 9808
rect 7314 9802 7320 9808
rect 11256 9802 11262 9808
rect 11314 9802 11320 9808
rect 15256 9802 15262 9808
rect 15314 9802 15320 9808
rect 19256 9802 19262 9808
rect 19314 9802 19320 9808
rect 23256 9802 23262 9808
rect 23314 9802 23320 9808
rect 27256 9802 27262 9808
rect 27314 9802 27320 9808
rect 31256 9802 31262 9808
rect 31314 9802 31320 9808
rect 35256 9802 35262 9808
rect 35314 9802 35320 9808
rect 39256 9802 39262 9808
rect 39314 9802 39320 9808
rect 3256 9756 3262 9762
rect 3314 9756 3320 9762
rect 7256 9756 7262 9762
rect 7314 9756 7320 9762
rect 11256 9756 11262 9762
rect 11314 9756 11320 9762
rect 15256 9756 15262 9762
rect 15314 9756 15320 9762
rect 19256 9756 19262 9762
rect 19314 9756 19320 9762
rect 23256 9756 23262 9762
rect 23314 9756 23320 9762
rect 27256 9756 27262 9762
rect 27314 9756 27320 9762
rect 31256 9756 31262 9762
rect 31314 9756 31320 9762
rect 35256 9756 35262 9762
rect 35314 9756 35320 9762
rect 39256 9756 39262 9762
rect 39314 9756 39320 9762
rect 3262 9750 3268 9756
rect 3308 9750 3314 9756
rect 7262 9750 7268 9756
rect 7308 9750 7314 9756
rect 11262 9750 11268 9756
rect 11308 9750 11314 9756
rect 15262 9750 15268 9756
rect 15308 9750 15314 9756
rect 19262 9750 19268 9756
rect 19308 9750 19314 9756
rect 23262 9750 23268 9756
rect 23308 9750 23314 9756
rect 27262 9750 27268 9756
rect 27308 9750 27314 9756
rect 31262 9750 31268 9756
rect 31308 9750 31314 9756
rect 35262 9750 35268 9756
rect 35308 9750 35314 9756
rect 39262 9750 39268 9756
rect 39308 9750 39314 9756
rect 2240 9296 2480 9320
rect 2240 9104 2264 9296
rect 2456 9104 2480 9296
rect 2240 9080 2480 9104
rect 6240 9296 6480 9320
rect 6240 9104 6264 9296
rect 6456 9104 6480 9296
rect 6240 9080 6480 9104
rect 10240 9296 10480 9320
rect 10240 9104 10264 9296
rect 10456 9104 10480 9296
rect 10240 9080 10480 9104
rect 14240 9296 14480 9320
rect 14240 9104 14264 9296
rect 14456 9104 14480 9296
rect 14240 9080 14480 9104
rect 18240 9296 18480 9320
rect 18240 9104 18264 9296
rect 18456 9104 18480 9296
rect 18240 9080 18480 9104
rect 22240 9296 22480 9320
rect 22240 9104 22264 9296
rect 22456 9104 22480 9296
rect 22240 9080 22480 9104
rect 26240 9296 26480 9320
rect 26240 9104 26264 9296
rect 26456 9104 26480 9296
rect 26240 9080 26480 9104
rect 30240 9296 30480 9320
rect 30240 9104 30264 9296
rect 30456 9104 30480 9296
rect 30240 9080 30480 9104
rect 34240 9296 34480 9320
rect 34240 9104 34264 9296
rect 34456 9104 34480 9296
rect 34240 9080 34480 9104
rect 38240 9296 38480 9320
rect 38240 9104 38264 9296
rect 38456 9104 38480 9296
rect 38240 9080 38480 9104
rect 2240 8596 2480 8620
rect 2240 8536 2264 8596
rect 2456 8536 2480 8596
rect 2240 8380 2480 8536
rect 6240 8596 6480 8620
rect 6240 8536 6264 8596
rect 6456 8536 6480 8596
rect 6240 8380 6480 8536
rect 10240 8596 10480 8620
rect 10240 8536 10264 8596
rect 10456 8536 10480 8596
rect 10240 8380 10480 8536
rect 14240 8596 14480 8620
rect 14240 8536 14264 8596
rect 14456 8536 14480 8596
rect 14240 8380 14480 8536
rect 18240 8596 18480 8620
rect 18240 8536 18264 8596
rect 18456 8536 18480 8596
rect 18240 8380 18480 8536
rect 22240 8596 22480 8620
rect 22240 8536 22264 8596
rect 22456 8536 22480 8596
rect 22240 8380 22480 8536
rect 26240 8596 26480 8620
rect 26240 8536 26264 8596
rect 26456 8536 26480 8596
rect 26240 8380 26480 8536
rect 30240 8596 30480 8620
rect 30240 8536 30264 8596
rect 30456 8536 30480 8596
rect 30240 8380 30480 8536
rect 34240 8596 34480 8620
rect 34240 8536 34264 8596
rect 34456 8536 34480 8596
rect 34240 8380 34480 8536
rect 38240 8596 38480 8620
rect 38240 8536 38264 8596
rect 38456 8536 38480 8596
rect 38240 8380 38480 8536
rect 1936 8160 2256 8216
rect 360 7916 600 7940
rect 360 7724 384 7916
rect 576 7724 600 7916
rect 1936 7920 1960 8160
rect 2224 7920 2256 8160
rect 3602 8163 3690 8168
rect 3602 8085 3607 8163
rect 3685 8085 3690 8163
rect 3602 8080 3690 8085
rect 5936 8160 6256 8216
rect 1936 7896 2256 7920
rect 4360 7916 4600 7940
rect 360 7700 600 7724
rect 4360 7724 4384 7916
rect 4576 7724 4600 7916
rect 5936 7920 5960 8160
rect 6224 7920 6256 8160
rect 7602 8163 7690 8168
rect 7602 8085 7607 8163
rect 7685 8085 7690 8163
rect 7602 8080 7690 8085
rect 9936 8160 10256 8216
rect 5936 7896 6256 7920
rect 8360 7916 8600 7940
rect 2810 7711 2946 7716
rect 2810 7637 2815 7711
rect 2941 7637 2946 7711
rect 4360 7700 4600 7724
rect 8360 7724 8384 7916
rect 8576 7724 8600 7916
rect 9936 7920 9960 8160
rect 10224 7920 10256 8160
rect 11602 8163 11690 8168
rect 11602 8085 11607 8163
rect 11685 8085 11690 8163
rect 11602 8080 11690 8085
rect 13936 8160 14256 8216
rect 9936 7896 10256 7920
rect 12360 7916 12600 7940
rect 6810 7711 6946 7716
rect 2810 7632 2946 7637
rect 6810 7637 6815 7711
rect 6941 7637 6946 7711
rect 8360 7700 8600 7724
rect 12360 7724 12384 7916
rect 12576 7724 12600 7916
rect 13936 7920 13960 8160
rect 14224 7920 14256 8160
rect 15602 8163 15690 8168
rect 15602 8085 15607 8163
rect 15685 8085 15690 8163
rect 15602 8080 15690 8085
rect 17936 8160 18256 8216
rect 13936 7896 14256 7920
rect 16360 7916 16600 7940
rect 10810 7711 10946 7716
rect 6810 7632 6946 7637
rect 10810 7637 10815 7711
rect 10941 7637 10946 7711
rect 12360 7700 12600 7724
rect 16360 7724 16384 7916
rect 16576 7724 16600 7916
rect 17936 7920 17960 8160
rect 18224 7920 18256 8160
rect 19602 8163 19690 8168
rect 19602 8085 19607 8163
rect 19685 8085 19690 8163
rect 19602 8080 19690 8085
rect 21936 8160 22256 8216
rect 17936 7896 18256 7920
rect 20360 7916 20600 7940
rect 14810 7711 14946 7716
rect 10810 7632 10946 7637
rect 14810 7637 14815 7711
rect 14941 7637 14946 7711
rect 16360 7700 16600 7724
rect 20360 7724 20384 7916
rect 20576 7724 20600 7916
rect 21936 7920 21960 8160
rect 22224 7920 22256 8160
rect 23602 8163 23690 8168
rect 23602 8085 23607 8163
rect 23685 8085 23690 8163
rect 23602 8080 23690 8085
rect 25936 8160 26256 8216
rect 21936 7896 22256 7920
rect 24360 7916 24600 7940
rect 18810 7711 18946 7716
rect 14810 7632 14946 7637
rect 18810 7637 18815 7711
rect 18941 7637 18946 7711
rect 20360 7700 20600 7724
rect 24360 7724 24384 7916
rect 24576 7724 24600 7916
rect 25936 7920 25960 8160
rect 26224 7920 26256 8160
rect 27602 8163 27690 8168
rect 27602 8085 27607 8163
rect 27685 8085 27690 8163
rect 27602 8080 27690 8085
rect 29936 8160 30256 8216
rect 25936 7896 26256 7920
rect 28360 7916 28600 7940
rect 22810 7711 22946 7716
rect 18810 7632 18946 7637
rect 22810 7637 22815 7711
rect 22941 7637 22946 7711
rect 24360 7700 24600 7724
rect 28360 7724 28384 7916
rect 28576 7724 28600 7916
rect 29936 7920 29960 8160
rect 30224 7920 30256 8160
rect 31602 8163 31690 8168
rect 31602 8085 31607 8163
rect 31685 8085 31690 8163
rect 31602 8080 31690 8085
rect 33936 8160 34256 8216
rect 29936 7896 30256 7920
rect 32360 7916 32600 7940
rect 26810 7711 26946 7716
rect 22810 7632 22946 7637
rect 26810 7637 26815 7711
rect 26941 7637 26946 7711
rect 28360 7700 28600 7724
rect 32360 7724 32384 7916
rect 32576 7724 32600 7916
rect 33936 7920 33960 8160
rect 34224 7920 34256 8160
rect 35602 8163 35690 8168
rect 35602 8085 35607 8163
rect 35685 8085 35690 8163
rect 35602 8080 35690 8085
rect 37936 8160 38256 8216
rect 33936 7896 34256 7920
rect 36360 7916 36600 7940
rect 30810 7711 30946 7716
rect 26810 7632 26946 7637
rect 30810 7637 30815 7711
rect 30941 7637 30946 7711
rect 32360 7700 32600 7724
rect 36360 7724 36384 7916
rect 36576 7724 36600 7916
rect 37936 7920 37960 8160
rect 38224 7920 38256 8160
rect 39602 8163 39690 8168
rect 39602 8085 39607 8163
rect 39685 8085 39690 8163
rect 39602 8080 39690 8085
rect 37936 7896 38256 7920
rect 34810 7711 34946 7716
rect 30810 7632 30946 7637
rect 34810 7637 34815 7711
rect 34941 7637 34946 7711
rect 36360 7700 36600 7724
rect 38810 7711 38946 7716
rect 34810 7632 34946 7637
rect 38810 7637 38815 7711
rect 38941 7637 38946 7711
rect 38810 7632 38946 7637
rect 2338 7573 2518 7574
rect 2338 7395 2339 7573
rect 2517 7395 2518 7573
rect 2338 7394 2518 7395
rect 6338 7573 6518 7574
rect 6338 7395 6339 7573
rect 6517 7395 6518 7573
rect 6338 7394 6518 7395
rect 10338 7573 10518 7574
rect 10338 7395 10339 7573
rect 10517 7395 10518 7573
rect 10338 7394 10518 7395
rect 14338 7573 14518 7574
rect 14338 7395 14339 7573
rect 14517 7395 14518 7573
rect 14338 7394 14518 7395
rect 18338 7573 18518 7574
rect 18338 7395 18339 7573
rect 18517 7395 18518 7573
rect 18338 7394 18518 7395
rect 22338 7573 22518 7574
rect 22338 7395 22339 7573
rect 22517 7395 22518 7573
rect 22338 7394 22518 7395
rect 26338 7573 26518 7574
rect 26338 7395 26339 7573
rect 26517 7395 26518 7573
rect 26338 7394 26518 7395
rect 30338 7573 30518 7574
rect 30338 7395 30339 7573
rect 30517 7395 30518 7573
rect 30338 7394 30518 7395
rect 34338 7573 34518 7574
rect 34338 7395 34339 7573
rect 34517 7395 34518 7573
rect 34338 7394 34518 7395
rect 38338 7573 38518 7574
rect 38338 7395 38339 7573
rect 38517 7395 38518 7573
rect 38338 7394 38518 7395
rect 400 6999 580 7000
rect 400 6821 401 6999
rect 579 6821 580 6999
rect 3734 6996 3740 7002
rect 3780 6996 3786 7002
rect 4400 6999 4580 7000
rect 3728 6990 3734 6996
rect 3786 6990 3792 6996
rect 3728 6944 3734 6950
rect 3786 6944 3792 6950
rect 3734 6938 3740 6944
rect 3780 6938 3786 6944
rect 400 6820 580 6821
rect 4400 6821 4401 6999
rect 4579 6821 4580 6999
rect 7734 6996 7740 7002
rect 7780 6996 7786 7002
rect 8400 6999 8580 7000
rect 7728 6990 7734 6996
rect 7786 6990 7792 6996
rect 7728 6944 7734 6950
rect 7786 6944 7792 6950
rect 7734 6938 7740 6944
rect 7780 6938 7786 6944
rect 4400 6820 4580 6821
rect 8400 6821 8401 6999
rect 8579 6821 8580 6999
rect 11734 6996 11740 7002
rect 11780 6996 11786 7002
rect 12400 6999 12580 7000
rect 11728 6990 11734 6996
rect 11786 6990 11792 6996
rect 11728 6944 11734 6950
rect 11786 6944 11792 6950
rect 11734 6938 11740 6944
rect 11780 6938 11786 6944
rect 8400 6820 8580 6821
rect 12400 6821 12401 6999
rect 12579 6821 12580 6999
rect 15734 6996 15740 7002
rect 15780 6996 15786 7002
rect 16400 6999 16580 7000
rect 15728 6990 15734 6996
rect 15786 6990 15792 6996
rect 15728 6944 15734 6950
rect 15786 6944 15792 6950
rect 15734 6938 15740 6944
rect 15780 6938 15786 6944
rect 12400 6820 12580 6821
rect 16400 6821 16401 6999
rect 16579 6821 16580 6999
rect 19734 6996 19740 7002
rect 19780 6996 19786 7002
rect 20400 6999 20580 7000
rect 19728 6990 19734 6996
rect 19786 6990 19792 6996
rect 19728 6944 19734 6950
rect 19786 6944 19792 6950
rect 19734 6938 19740 6944
rect 19780 6938 19786 6944
rect 16400 6820 16580 6821
rect 20400 6821 20401 6999
rect 20579 6821 20580 6999
rect 23734 6996 23740 7002
rect 23780 6996 23786 7002
rect 24400 6999 24580 7000
rect 23728 6990 23734 6996
rect 23786 6990 23792 6996
rect 23728 6944 23734 6950
rect 23786 6944 23792 6950
rect 23734 6938 23740 6944
rect 23780 6938 23786 6944
rect 20400 6820 20580 6821
rect 24400 6821 24401 6999
rect 24579 6821 24580 6999
rect 27734 6996 27740 7002
rect 27780 6996 27786 7002
rect 28400 6999 28580 7000
rect 27728 6990 27734 6996
rect 27786 6990 27792 6996
rect 27728 6944 27734 6950
rect 27786 6944 27792 6950
rect 27734 6938 27740 6944
rect 27780 6938 27786 6944
rect 24400 6820 24580 6821
rect 28400 6821 28401 6999
rect 28579 6821 28580 6999
rect 31734 6996 31740 7002
rect 31780 6996 31786 7002
rect 32400 6999 32580 7000
rect 31728 6990 31734 6996
rect 31786 6990 31792 6996
rect 31728 6944 31734 6950
rect 31786 6944 31792 6950
rect 31734 6938 31740 6944
rect 31780 6938 31786 6944
rect 28400 6820 28580 6821
rect 32400 6821 32401 6999
rect 32579 6821 32580 6999
rect 35734 6996 35740 7002
rect 35780 6996 35786 7002
rect 36400 6999 36580 7000
rect 35728 6990 35734 6996
rect 35786 6990 35792 6996
rect 35728 6944 35734 6950
rect 35786 6944 35792 6950
rect 35734 6938 35740 6944
rect 35780 6938 35786 6944
rect 32400 6820 32580 6821
rect 36400 6821 36401 6999
rect 36579 6821 36580 6999
rect 39734 6996 39740 7002
rect 39780 6996 39786 7002
rect 39728 6990 39734 6996
rect 39786 6990 39792 6996
rect 39728 6944 39734 6950
rect 39786 6944 39792 6950
rect 39734 6938 39740 6944
rect 39780 6938 39786 6944
rect 36400 6820 36580 6821
rect 3262 6808 3268 6814
rect 3308 6808 3314 6814
rect 7262 6808 7268 6814
rect 7308 6808 7314 6814
rect 11262 6808 11268 6814
rect 11308 6808 11314 6814
rect 15262 6808 15268 6814
rect 15308 6808 15314 6814
rect 19262 6808 19268 6814
rect 19308 6808 19314 6814
rect 23262 6808 23268 6814
rect 23308 6808 23314 6814
rect 27262 6808 27268 6814
rect 27308 6808 27314 6814
rect 31262 6808 31268 6814
rect 31308 6808 31314 6814
rect 35262 6808 35268 6814
rect 35308 6808 35314 6814
rect 39262 6808 39268 6814
rect 39308 6808 39314 6814
rect 3256 6802 3262 6808
rect 3314 6802 3320 6808
rect 7256 6802 7262 6808
rect 7314 6802 7320 6808
rect 11256 6802 11262 6808
rect 11314 6802 11320 6808
rect 15256 6802 15262 6808
rect 15314 6802 15320 6808
rect 19256 6802 19262 6808
rect 19314 6802 19320 6808
rect 23256 6802 23262 6808
rect 23314 6802 23320 6808
rect 27256 6802 27262 6808
rect 27314 6802 27320 6808
rect 31256 6802 31262 6808
rect 31314 6802 31320 6808
rect 35256 6802 35262 6808
rect 35314 6802 35320 6808
rect 39256 6802 39262 6808
rect 39314 6802 39320 6808
rect 3256 6756 3262 6762
rect 3314 6756 3320 6762
rect 7256 6756 7262 6762
rect 7314 6756 7320 6762
rect 11256 6756 11262 6762
rect 11314 6756 11320 6762
rect 15256 6756 15262 6762
rect 15314 6756 15320 6762
rect 19256 6756 19262 6762
rect 19314 6756 19320 6762
rect 23256 6756 23262 6762
rect 23314 6756 23320 6762
rect 27256 6756 27262 6762
rect 27314 6756 27320 6762
rect 31256 6756 31262 6762
rect 31314 6756 31320 6762
rect 35256 6756 35262 6762
rect 35314 6756 35320 6762
rect 39256 6756 39262 6762
rect 39314 6756 39320 6762
rect 3262 6750 3268 6756
rect 3308 6750 3314 6756
rect 7262 6750 7268 6756
rect 7308 6750 7314 6756
rect 11262 6750 11268 6756
rect 11308 6750 11314 6756
rect 15262 6750 15268 6756
rect 15308 6750 15314 6756
rect 19262 6750 19268 6756
rect 19308 6750 19314 6756
rect 23262 6750 23268 6756
rect 23308 6750 23314 6756
rect 27262 6750 27268 6756
rect 27308 6750 27314 6756
rect 31262 6750 31268 6756
rect 31308 6750 31314 6756
rect 35262 6750 35268 6756
rect 35308 6750 35314 6756
rect 39262 6750 39268 6756
rect 39308 6750 39314 6756
rect 2240 6296 2480 6320
rect 2240 6104 2264 6296
rect 2456 6104 2480 6296
rect 2240 6080 2480 6104
rect 6240 6296 6480 6320
rect 6240 6104 6264 6296
rect 6456 6104 6480 6296
rect 6240 6080 6480 6104
rect 10240 6296 10480 6320
rect 10240 6104 10264 6296
rect 10456 6104 10480 6296
rect 10240 6080 10480 6104
rect 14240 6296 14480 6320
rect 14240 6104 14264 6296
rect 14456 6104 14480 6296
rect 14240 6080 14480 6104
rect 18240 6296 18480 6320
rect 18240 6104 18264 6296
rect 18456 6104 18480 6296
rect 18240 6080 18480 6104
rect 22240 6296 22480 6320
rect 22240 6104 22264 6296
rect 22456 6104 22480 6296
rect 22240 6080 22480 6104
rect 26240 6296 26480 6320
rect 26240 6104 26264 6296
rect 26456 6104 26480 6296
rect 26240 6080 26480 6104
rect 30240 6296 30480 6320
rect 30240 6104 30264 6296
rect 30456 6104 30480 6296
rect 30240 6080 30480 6104
rect 34240 6296 34480 6320
rect 34240 6104 34264 6296
rect 34456 6104 34480 6296
rect 34240 6080 34480 6104
rect 38240 6296 38480 6320
rect 38240 6104 38264 6296
rect 38456 6104 38480 6296
rect 38240 6080 38480 6104
rect 2240 5596 2480 5620
rect 2240 5536 2264 5596
rect 2456 5536 2480 5596
rect 2240 5380 2480 5536
rect 6240 5596 6480 5620
rect 6240 5536 6264 5596
rect 6456 5536 6480 5596
rect 6240 5380 6480 5536
rect 10240 5596 10480 5620
rect 10240 5536 10264 5596
rect 10456 5536 10480 5596
rect 10240 5380 10480 5536
rect 14240 5596 14480 5620
rect 14240 5536 14264 5596
rect 14456 5536 14480 5596
rect 14240 5380 14480 5536
rect 18240 5596 18480 5620
rect 18240 5536 18264 5596
rect 18456 5536 18480 5596
rect 18240 5380 18480 5536
rect 22240 5596 22480 5620
rect 22240 5536 22264 5596
rect 22456 5536 22480 5596
rect 22240 5380 22480 5536
rect 26240 5596 26480 5620
rect 26240 5536 26264 5596
rect 26456 5536 26480 5596
rect 26240 5380 26480 5536
rect 30240 5596 30480 5620
rect 30240 5536 30264 5596
rect 30456 5536 30480 5596
rect 30240 5380 30480 5536
rect 34240 5596 34480 5620
rect 34240 5536 34264 5596
rect 34456 5536 34480 5596
rect 34240 5380 34480 5536
rect 38240 5596 38480 5620
rect 38240 5536 38264 5596
rect 38456 5536 38480 5596
rect 38240 5380 38480 5536
rect 1936 5160 2256 5216
rect 360 4916 600 4940
rect 360 4724 384 4916
rect 576 4724 600 4916
rect 1936 4920 1960 5160
rect 2224 4920 2256 5160
rect 3602 5163 3690 5168
rect 3602 5085 3607 5163
rect 3685 5085 3690 5163
rect 3602 5080 3690 5085
rect 5936 5160 6256 5216
rect 1936 4896 2256 4920
rect 4360 4916 4600 4940
rect 360 4700 600 4724
rect 4360 4724 4384 4916
rect 4576 4724 4600 4916
rect 5936 4920 5960 5160
rect 6224 4920 6256 5160
rect 7602 5163 7690 5168
rect 7602 5085 7607 5163
rect 7685 5085 7690 5163
rect 7602 5080 7690 5085
rect 9936 5160 10256 5216
rect 5936 4896 6256 4920
rect 8360 4916 8600 4940
rect 2810 4711 2946 4716
rect 2810 4637 2815 4711
rect 2941 4637 2946 4711
rect 4360 4700 4600 4724
rect 8360 4724 8384 4916
rect 8576 4724 8600 4916
rect 9936 4920 9960 5160
rect 10224 4920 10256 5160
rect 11602 5163 11690 5168
rect 11602 5085 11607 5163
rect 11685 5085 11690 5163
rect 11602 5080 11690 5085
rect 13936 5160 14256 5216
rect 9936 4896 10256 4920
rect 12360 4916 12600 4940
rect 6810 4711 6946 4716
rect 2810 4632 2946 4637
rect 6810 4637 6815 4711
rect 6941 4637 6946 4711
rect 8360 4700 8600 4724
rect 12360 4724 12384 4916
rect 12576 4724 12600 4916
rect 13936 4920 13960 5160
rect 14224 4920 14256 5160
rect 15602 5163 15690 5168
rect 15602 5085 15607 5163
rect 15685 5085 15690 5163
rect 15602 5080 15690 5085
rect 17936 5160 18256 5216
rect 13936 4896 14256 4920
rect 16360 4916 16600 4940
rect 10810 4711 10946 4716
rect 6810 4632 6946 4637
rect 10810 4637 10815 4711
rect 10941 4637 10946 4711
rect 12360 4700 12600 4724
rect 16360 4724 16384 4916
rect 16576 4724 16600 4916
rect 17936 4920 17960 5160
rect 18224 4920 18256 5160
rect 19602 5163 19690 5168
rect 19602 5085 19607 5163
rect 19685 5085 19690 5163
rect 19602 5080 19690 5085
rect 21936 5160 22256 5216
rect 17936 4896 18256 4920
rect 20360 4916 20600 4940
rect 14810 4711 14946 4716
rect 10810 4632 10946 4637
rect 14810 4637 14815 4711
rect 14941 4637 14946 4711
rect 16360 4700 16600 4724
rect 20360 4724 20384 4916
rect 20576 4724 20600 4916
rect 21936 4920 21960 5160
rect 22224 4920 22256 5160
rect 23602 5163 23690 5168
rect 23602 5085 23607 5163
rect 23685 5085 23690 5163
rect 23602 5080 23690 5085
rect 25936 5160 26256 5216
rect 21936 4896 22256 4920
rect 24360 4916 24600 4940
rect 18810 4711 18946 4716
rect 14810 4632 14946 4637
rect 18810 4637 18815 4711
rect 18941 4637 18946 4711
rect 20360 4700 20600 4724
rect 24360 4724 24384 4916
rect 24576 4724 24600 4916
rect 25936 4920 25960 5160
rect 26224 4920 26256 5160
rect 27602 5163 27690 5168
rect 27602 5085 27607 5163
rect 27685 5085 27690 5163
rect 27602 5080 27690 5085
rect 29936 5160 30256 5216
rect 25936 4896 26256 4920
rect 28360 4916 28600 4940
rect 22810 4711 22946 4716
rect 18810 4632 18946 4637
rect 22810 4637 22815 4711
rect 22941 4637 22946 4711
rect 24360 4700 24600 4724
rect 28360 4724 28384 4916
rect 28576 4724 28600 4916
rect 29936 4920 29960 5160
rect 30224 4920 30256 5160
rect 31602 5163 31690 5168
rect 31602 5085 31607 5163
rect 31685 5085 31690 5163
rect 31602 5080 31690 5085
rect 33936 5160 34256 5216
rect 29936 4896 30256 4920
rect 32360 4916 32600 4940
rect 26810 4711 26946 4716
rect 22810 4632 22946 4637
rect 26810 4637 26815 4711
rect 26941 4637 26946 4711
rect 28360 4700 28600 4724
rect 32360 4724 32384 4916
rect 32576 4724 32600 4916
rect 33936 4920 33960 5160
rect 34224 4920 34256 5160
rect 35602 5163 35690 5168
rect 35602 5085 35607 5163
rect 35685 5085 35690 5163
rect 35602 5080 35690 5085
rect 37936 5160 38256 5216
rect 33936 4896 34256 4920
rect 36360 4916 36600 4940
rect 30810 4711 30946 4716
rect 26810 4632 26946 4637
rect 30810 4637 30815 4711
rect 30941 4637 30946 4711
rect 32360 4700 32600 4724
rect 36360 4724 36384 4916
rect 36576 4724 36600 4916
rect 37936 4920 37960 5160
rect 38224 4920 38256 5160
rect 39602 5163 39690 5168
rect 39602 5085 39607 5163
rect 39685 5085 39690 5163
rect 39602 5080 39690 5085
rect 37936 4896 38256 4920
rect 34810 4711 34946 4716
rect 30810 4632 30946 4637
rect 34810 4637 34815 4711
rect 34941 4637 34946 4711
rect 36360 4700 36600 4724
rect 38810 4711 38946 4716
rect 34810 4632 34946 4637
rect 38810 4637 38815 4711
rect 38941 4637 38946 4711
rect 38810 4632 38946 4637
rect 2338 4573 2518 4574
rect 2338 4395 2339 4573
rect 2517 4395 2518 4573
rect 2338 4394 2518 4395
rect 6338 4573 6518 4574
rect 6338 4395 6339 4573
rect 6517 4395 6518 4573
rect 6338 4394 6518 4395
rect 10338 4573 10518 4574
rect 10338 4395 10339 4573
rect 10517 4395 10518 4573
rect 10338 4394 10518 4395
rect 14338 4573 14518 4574
rect 14338 4395 14339 4573
rect 14517 4395 14518 4573
rect 14338 4394 14518 4395
rect 18338 4573 18518 4574
rect 18338 4395 18339 4573
rect 18517 4395 18518 4573
rect 18338 4394 18518 4395
rect 22338 4573 22518 4574
rect 22338 4395 22339 4573
rect 22517 4395 22518 4573
rect 22338 4394 22518 4395
rect 26338 4573 26518 4574
rect 26338 4395 26339 4573
rect 26517 4395 26518 4573
rect 26338 4394 26518 4395
rect 30338 4573 30518 4574
rect 30338 4395 30339 4573
rect 30517 4395 30518 4573
rect 30338 4394 30518 4395
rect 34338 4573 34518 4574
rect 34338 4395 34339 4573
rect 34517 4395 34518 4573
rect 34338 4394 34518 4395
rect 38338 4573 38518 4574
rect 38338 4395 38339 4573
rect 38517 4395 38518 4573
rect 38338 4394 38518 4395
rect 400 3999 580 4000
rect 400 3821 401 3999
rect 579 3821 580 3999
rect 3734 3996 3740 4002
rect 3780 3996 3786 4002
rect 4400 3999 4580 4000
rect 3728 3990 3734 3996
rect 3786 3990 3792 3996
rect 3728 3944 3734 3950
rect 3786 3944 3792 3950
rect 3734 3938 3740 3944
rect 3780 3938 3786 3944
rect 400 3820 580 3821
rect 4400 3821 4401 3999
rect 4579 3821 4580 3999
rect 7734 3996 7740 4002
rect 7780 3996 7786 4002
rect 8400 3999 8580 4000
rect 7728 3990 7734 3996
rect 7786 3990 7792 3996
rect 7728 3944 7734 3950
rect 7786 3944 7792 3950
rect 7734 3938 7740 3944
rect 7780 3938 7786 3944
rect 4400 3820 4580 3821
rect 8400 3821 8401 3999
rect 8579 3821 8580 3999
rect 11734 3996 11740 4002
rect 11780 3996 11786 4002
rect 12400 3999 12580 4000
rect 11728 3990 11734 3996
rect 11786 3990 11792 3996
rect 11728 3944 11734 3950
rect 11786 3944 11792 3950
rect 11734 3938 11740 3944
rect 11780 3938 11786 3944
rect 8400 3820 8580 3821
rect 12400 3821 12401 3999
rect 12579 3821 12580 3999
rect 15734 3996 15740 4002
rect 15780 3996 15786 4002
rect 16400 3999 16580 4000
rect 15728 3990 15734 3996
rect 15786 3990 15792 3996
rect 15728 3944 15734 3950
rect 15786 3944 15792 3950
rect 15734 3938 15740 3944
rect 15780 3938 15786 3944
rect 12400 3820 12580 3821
rect 16400 3821 16401 3999
rect 16579 3821 16580 3999
rect 19734 3996 19740 4002
rect 19780 3996 19786 4002
rect 20400 3999 20580 4000
rect 19728 3990 19734 3996
rect 19786 3990 19792 3996
rect 19728 3944 19734 3950
rect 19786 3944 19792 3950
rect 19734 3938 19740 3944
rect 19780 3938 19786 3944
rect 16400 3820 16580 3821
rect 20400 3821 20401 3999
rect 20579 3821 20580 3999
rect 23734 3996 23740 4002
rect 23780 3996 23786 4002
rect 24400 3999 24580 4000
rect 23728 3990 23734 3996
rect 23786 3990 23792 3996
rect 23728 3944 23734 3950
rect 23786 3944 23792 3950
rect 23734 3938 23740 3944
rect 23780 3938 23786 3944
rect 20400 3820 20580 3821
rect 24400 3821 24401 3999
rect 24579 3821 24580 3999
rect 27734 3996 27740 4002
rect 27780 3996 27786 4002
rect 28400 3999 28580 4000
rect 27728 3990 27734 3996
rect 27786 3990 27792 3996
rect 27728 3944 27734 3950
rect 27786 3944 27792 3950
rect 27734 3938 27740 3944
rect 27780 3938 27786 3944
rect 24400 3820 24580 3821
rect 28400 3821 28401 3999
rect 28579 3821 28580 3999
rect 31734 3996 31740 4002
rect 31780 3996 31786 4002
rect 32400 3999 32580 4000
rect 31728 3990 31734 3996
rect 31786 3990 31792 3996
rect 31728 3944 31734 3950
rect 31786 3944 31792 3950
rect 31734 3938 31740 3944
rect 31780 3938 31786 3944
rect 28400 3820 28580 3821
rect 32400 3821 32401 3999
rect 32579 3821 32580 3999
rect 35734 3996 35740 4002
rect 35780 3996 35786 4002
rect 36400 3999 36580 4000
rect 35728 3990 35734 3996
rect 35786 3990 35792 3996
rect 35728 3944 35734 3950
rect 35786 3944 35792 3950
rect 35734 3938 35740 3944
rect 35780 3938 35786 3944
rect 32400 3820 32580 3821
rect 36400 3821 36401 3999
rect 36579 3821 36580 3999
rect 39734 3996 39740 4002
rect 39780 3996 39786 4002
rect 39728 3990 39734 3996
rect 39786 3990 39792 3996
rect 39728 3944 39734 3950
rect 39786 3944 39792 3950
rect 39734 3938 39740 3944
rect 39780 3938 39786 3944
rect 36400 3820 36580 3821
rect 3262 3808 3268 3814
rect 3308 3808 3314 3814
rect 7262 3808 7268 3814
rect 7308 3808 7314 3814
rect 11262 3808 11268 3814
rect 11308 3808 11314 3814
rect 15262 3808 15268 3814
rect 15308 3808 15314 3814
rect 19262 3808 19268 3814
rect 19308 3808 19314 3814
rect 23262 3808 23268 3814
rect 23308 3808 23314 3814
rect 27262 3808 27268 3814
rect 27308 3808 27314 3814
rect 31262 3808 31268 3814
rect 31308 3808 31314 3814
rect 35262 3808 35268 3814
rect 35308 3808 35314 3814
rect 39262 3808 39268 3814
rect 39308 3808 39314 3814
rect 3256 3802 3262 3808
rect 3314 3802 3320 3808
rect 7256 3802 7262 3808
rect 7314 3802 7320 3808
rect 11256 3802 11262 3808
rect 11314 3802 11320 3808
rect 15256 3802 15262 3808
rect 15314 3802 15320 3808
rect 19256 3802 19262 3808
rect 19314 3802 19320 3808
rect 23256 3802 23262 3808
rect 23314 3802 23320 3808
rect 27256 3802 27262 3808
rect 27314 3802 27320 3808
rect 31256 3802 31262 3808
rect 31314 3802 31320 3808
rect 35256 3802 35262 3808
rect 35314 3802 35320 3808
rect 39256 3802 39262 3808
rect 39314 3802 39320 3808
rect 3256 3756 3262 3762
rect 3314 3756 3320 3762
rect 7256 3756 7262 3762
rect 7314 3756 7320 3762
rect 11256 3756 11262 3762
rect 11314 3756 11320 3762
rect 15256 3756 15262 3762
rect 15314 3756 15320 3762
rect 19256 3756 19262 3762
rect 19314 3756 19320 3762
rect 23256 3756 23262 3762
rect 23314 3756 23320 3762
rect 27256 3756 27262 3762
rect 27314 3756 27320 3762
rect 31256 3756 31262 3762
rect 31314 3756 31320 3762
rect 35256 3756 35262 3762
rect 35314 3756 35320 3762
rect 39256 3756 39262 3762
rect 39314 3756 39320 3762
rect 3262 3750 3268 3756
rect 3308 3750 3314 3756
rect 7262 3750 7268 3756
rect 7308 3750 7314 3756
rect 11262 3750 11268 3756
rect 11308 3750 11314 3756
rect 15262 3750 15268 3756
rect 15308 3750 15314 3756
rect 19262 3750 19268 3756
rect 19308 3750 19314 3756
rect 23262 3750 23268 3756
rect 23308 3750 23314 3756
rect 27262 3750 27268 3756
rect 27308 3750 27314 3756
rect 31262 3750 31268 3756
rect 31308 3750 31314 3756
rect 35262 3750 35268 3756
rect 35308 3750 35314 3756
rect 39262 3750 39268 3756
rect 39308 3750 39314 3756
rect 2240 3296 2480 3320
rect 2240 3104 2264 3296
rect 2456 3104 2480 3296
rect 2240 3080 2480 3104
rect 6240 3296 6480 3320
rect 6240 3104 6264 3296
rect 6456 3104 6480 3296
rect 6240 3080 6480 3104
rect 10240 3296 10480 3320
rect 10240 3104 10264 3296
rect 10456 3104 10480 3296
rect 10240 3080 10480 3104
rect 14240 3296 14480 3320
rect 14240 3104 14264 3296
rect 14456 3104 14480 3296
rect 14240 3080 14480 3104
rect 18240 3296 18480 3320
rect 18240 3104 18264 3296
rect 18456 3104 18480 3296
rect 18240 3080 18480 3104
rect 22240 3296 22480 3320
rect 22240 3104 22264 3296
rect 22456 3104 22480 3296
rect 22240 3080 22480 3104
rect 26240 3296 26480 3320
rect 26240 3104 26264 3296
rect 26456 3104 26480 3296
rect 26240 3080 26480 3104
rect 30240 3296 30480 3320
rect 30240 3104 30264 3296
rect 30456 3104 30480 3296
rect 30240 3080 30480 3104
rect 34240 3296 34480 3320
rect 34240 3104 34264 3296
rect 34456 3104 34480 3296
rect 34240 3080 34480 3104
rect 38240 3296 38480 3320
rect 38240 3104 38264 3296
rect 38456 3104 38480 3296
rect 38240 3080 38480 3104
rect 2240 2596 2480 2620
rect 2240 2536 2264 2596
rect 2456 2536 2480 2596
rect 2240 2380 2480 2536
rect 6240 2596 6480 2620
rect 6240 2536 6264 2596
rect 6456 2536 6480 2596
rect 6240 2380 6480 2536
rect 10240 2596 10480 2620
rect 10240 2536 10264 2596
rect 10456 2536 10480 2596
rect 10240 2380 10480 2536
rect 14240 2596 14480 2620
rect 14240 2536 14264 2596
rect 14456 2536 14480 2596
rect 14240 2380 14480 2536
rect 18240 2596 18480 2620
rect 18240 2536 18264 2596
rect 18456 2536 18480 2596
rect 18240 2380 18480 2536
rect 22240 2596 22480 2620
rect 22240 2536 22264 2596
rect 22456 2536 22480 2596
rect 22240 2380 22480 2536
rect 26240 2596 26480 2620
rect 26240 2536 26264 2596
rect 26456 2536 26480 2596
rect 26240 2380 26480 2536
rect 30240 2596 30480 2620
rect 30240 2536 30264 2596
rect 30456 2536 30480 2596
rect 30240 2380 30480 2536
rect 34240 2596 34480 2620
rect 34240 2536 34264 2596
rect 34456 2536 34480 2596
rect 34240 2380 34480 2536
rect 38240 2596 38480 2620
rect 38240 2536 38264 2596
rect 38456 2536 38480 2596
rect 38240 2380 38480 2536
rect 1936 2160 2256 2216
rect 360 1916 600 1940
rect 360 1724 384 1916
rect 576 1724 600 1916
rect 1936 1920 1960 2160
rect 2224 1920 2256 2160
rect 3602 2163 3690 2168
rect 3602 2085 3607 2163
rect 3685 2085 3690 2163
rect 3602 2080 3690 2085
rect 5936 2160 6256 2216
rect 1936 1896 2256 1920
rect 4360 1916 4600 1940
rect 360 1700 600 1724
rect 4360 1724 4384 1916
rect 4576 1724 4600 1916
rect 5936 1920 5960 2160
rect 6224 1920 6256 2160
rect 7602 2163 7690 2168
rect 7602 2085 7607 2163
rect 7685 2085 7690 2163
rect 7602 2080 7690 2085
rect 9936 2160 10256 2216
rect 5936 1896 6256 1920
rect 8360 1916 8600 1940
rect 2810 1711 2946 1716
rect 2810 1637 2815 1711
rect 2941 1637 2946 1711
rect 4360 1700 4600 1724
rect 8360 1724 8384 1916
rect 8576 1724 8600 1916
rect 9936 1920 9960 2160
rect 10224 1920 10256 2160
rect 11602 2163 11690 2168
rect 11602 2085 11607 2163
rect 11685 2085 11690 2163
rect 11602 2080 11690 2085
rect 13936 2160 14256 2216
rect 9936 1896 10256 1920
rect 12360 1916 12600 1940
rect 6810 1711 6946 1716
rect 2810 1632 2946 1637
rect 6810 1637 6815 1711
rect 6941 1637 6946 1711
rect 8360 1700 8600 1724
rect 12360 1724 12384 1916
rect 12576 1724 12600 1916
rect 13936 1920 13960 2160
rect 14224 1920 14256 2160
rect 15602 2163 15690 2168
rect 15602 2085 15607 2163
rect 15685 2085 15690 2163
rect 15602 2080 15690 2085
rect 17936 2160 18256 2216
rect 13936 1896 14256 1920
rect 16360 1916 16600 1940
rect 10810 1711 10946 1716
rect 6810 1632 6946 1637
rect 10810 1637 10815 1711
rect 10941 1637 10946 1711
rect 12360 1700 12600 1724
rect 16360 1724 16384 1916
rect 16576 1724 16600 1916
rect 17936 1920 17960 2160
rect 18224 1920 18256 2160
rect 19602 2163 19690 2168
rect 19602 2085 19607 2163
rect 19685 2085 19690 2163
rect 19602 2080 19690 2085
rect 21936 2160 22256 2216
rect 17936 1896 18256 1920
rect 20360 1916 20600 1940
rect 14810 1711 14946 1716
rect 10810 1632 10946 1637
rect 14810 1637 14815 1711
rect 14941 1637 14946 1711
rect 16360 1700 16600 1724
rect 20360 1724 20384 1916
rect 20576 1724 20600 1916
rect 21936 1920 21960 2160
rect 22224 1920 22256 2160
rect 23602 2163 23690 2168
rect 23602 2085 23607 2163
rect 23685 2085 23690 2163
rect 23602 2080 23690 2085
rect 25936 2160 26256 2216
rect 21936 1896 22256 1920
rect 24360 1916 24600 1940
rect 18810 1711 18946 1716
rect 14810 1632 14946 1637
rect 18810 1637 18815 1711
rect 18941 1637 18946 1711
rect 20360 1700 20600 1724
rect 24360 1724 24384 1916
rect 24576 1724 24600 1916
rect 25936 1920 25960 2160
rect 26224 1920 26256 2160
rect 27602 2163 27690 2168
rect 27602 2085 27607 2163
rect 27685 2085 27690 2163
rect 27602 2080 27690 2085
rect 29936 2160 30256 2216
rect 25936 1896 26256 1920
rect 28360 1916 28600 1940
rect 22810 1711 22946 1716
rect 18810 1632 18946 1637
rect 22810 1637 22815 1711
rect 22941 1637 22946 1711
rect 24360 1700 24600 1724
rect 28360 1724 28384 1916
rect 28576 1724 28600 1916
rect 29936 1920 29960 2160
rect 30224 1920 30256 2160
rect 31602 2163 31690 2168
rect 31602 2085 31607 2163
rect 31685 2085 31690 2163
rect 31602 2080 31690 2085
rect 33936 2160 34256 2216
rect 29936 1896 30256 1920
rect 32360 1916 32600 1940
rect 26810 1711 26946 1716
rect 22810 1632 22946 1637
rect 26810 1637 26815 1711
rect 26941 1637 26946 1711
rect 28360 1700 28600 1724
rect 32360 1724 32384 1916
rect 32576 1724 32600 1916
rect 33936 1920 33960 2160
rect 34224 1920 34256 2160
rect 35602 2163 35690 2168
rect 35602 2085 35607 2163
rect 35685 2085 35690 2163
rect 35602 2080 35690 2085
rect 37936 2160 38256 2216
rect 33936 1896 34256 1920
rect 36360 1916 36600 1940
rect 30810 1711 30946 1716
rect 26810 1632 26946 1637
rect 30810 1637 30815 1711
rect 30941 1637 30946 1711
rect 32360 1700 32600 1724
rect 36360 1724 36384 1916
rect 36576 1724 36600 1916
rect 37936 1920 37960 2160
rect 38224 1920 38256 2160
rect 39602 2163 39690 2168
rect 39602 2085 39607 2163
rect 39685 2085 39690 2163
rect 39602 2080 39690 2085
rect 37936 1896 38256 1920
rect 34810 1711 34946 1716
rect 30810 1632 30946 1637
rect 34810 1637 34815 1711
rect 34941 1637 34946 1711
rect 36360 1700 36600 1724
rect 38810 1711 38946 1716
rect 34810 1632 34946 1637
rect 38810 1637 38815 1711
rect 38941 1637 38946 1711
rect 38810 1632 38946 1637
rect 2338 1573 2518 1574
rect 2338 1395 2339 1573
rect 2517 1395 2518 1573
rect 2338 1394 2518 1395
rect 6338 1573 6518 1574
rect 6338 1395 6339 1573
rect 6517 1395 6518 1573
rect 6338 1394 6518 1395
rect 10338 1573 10518 1574
rect 10338 1395 10339 1573
rect 10517 1395 10518 1573
rect 10338 1394 10518 1395
rect 14338 1573 14518 1574
rect 14338 1395 14339 1573
rect 14517 1395 14518 1573
rect 14338 1394 14518 1395
rect 18338 1573 18518 1574
rect 18338 1395 18339 1573
rect 18517 1395 18518 1573
rect 18338 1394 18518 1395
rect 22338 1573 22518 1574
rect 22338 1395 22339 1573
rect 22517 1395 22518 1573
rect 22338 1394 22518 1395
rect 26338 1573 26518 1574
rect 26338 1395 26339 1573
rect 26517 1395 26518 1573
rect 26338 1394 26518 1395
rect 30338 1573 30518 1574
rect 30338 1395 30339 1573
rect 30517 1395 30518 1573
rect 30338 1394 30518 1395
rect 34338 1573 34518 1574
rect 34338 1395 34339 1573
rect 34517 1395 34518 1573
rect 34338 1394 34518 1395
rect 38338 1573 38518 1574
rect 38338 1395 38339 1573
rect 38517 1395 38518 1573
rect 38338 1394 38518 1395
rect 400 999 580 1000
rect 400 821 401 999
rect 579 821 580 999
rect 3734 996 3740 1002
rect 3780 996 3786 1002
rect 4400 999 4580 1000
rect 3728 990 3734 996
rect 3786 990 3792 996
rect 3728 944 3734 950
rect 3786 944 3792 950
rect 3734 938 3740 944
rect 3780 938 3786 944
rect 400 820 580 821
rect 4400 821 4401 999
rect 4579 821 4580 999
rect 7734 996 7740 1002
rect 7780 996 7786 1002
rect 8400 999 8580 1000
rect 7728 990 7734 996
rect 7786 990 7792 996
rect 7728 944 7734 950
rect 7786 944 7792 950
rect 7734 938 7740 944
rect 7780 938 7786 944
rect 4400 820 4580 821
rect 8400 821 8401 999
rect 8579 821 8580 999
rect 11734 996 11740 1002
rect 11780 996 11786 1002
rect 12400 999 12580 1000
rect 11728 990 11734 996
rect 11786 990 11792 996
rect 11728 944 11734 950
rect 11786 944 11792 950
rect 11734 938 11740 944
rect 11780 938 11786 944
rect 8400 820 8580 821
rect 12400 821 12401 999
rect 12579 821 12580 999
rect 15734 996 15740 1002
rect 15780 996 15786 1002
rect 16400 999 16580 1000
rect 15728 990 15734 996
rect 15786 990 15792 996
rect 15728 944 15734 950
rect 15786 944 15792 950
rect 15734 938 15740 944
rect 15780 938 15786 944
rect 12400 820 12580 821
rect 16400 821 16401 999
rect 16579 821 16580 999
rect 19734 996 19740 1002
rect 19780 996 19786 1002
rect 20400 999 20580 1000
rect 19728 990 19734 996
rect 19786 990 19792 996
rect 19728 944 19734 950
rect 19786 944 19792 950
rect 19734 938 19740 944
rect 19780 938 19786 944
rect 16400 820 16580 821
rect 20400 821 20401 999
rect 20579 821 20580 999
rect 23734 996 23740 1002
rect 23780 996 23786 1002
rect 24400 999 24580 1000
rect 23728 990 23734 996
rect 23786 990 23792 996
rect 23728 944 23734 950
rect 23786 944 23792 950
rect 23734 938 23740 944
rect 23780 938 23786 944
rect 20400 820 20580 821
rect 24400 821 24401 999
rect 24579 821 24580 999
rect 27734 996 27740 1002
rect 27780 996 27786 1002
rect 28400 999 28580 1000
rect 27728 990 27734 996
rect 27786 990 27792 996
rect 27728 944 27734 950
rect 27786 944 27792 950
rect 27734 938 27740 944
rect 27780 938 27786 944
rect 24400 820 24580 821
rect 28400 821 28401 999
rect 28579 821 28580 999
rect 31734 996 31740 1002
rect 31780 996 31786 1002
rect 32400 999 32580 1000
rect 31728 990 31734 996
rect 31786 990 31792 996
rect 31728 944 31734 950
rect 31786 944 31792 950
rect 31734 938 31740 944
rect 31780 938 31786 944
rect 28400 820 28580 821
rect 32400 821 32401 999
rect 32579 821 32580 999
rect 35734 996 35740 1002
rect 35780 996 35786 1002
rect 36400 999 36580 1000
rect 35728 990 35734 996
rect 35786 990 35792 996
rect 35728 944 35734 950
rect 35786 944 35792 950
rect 35734 938 35740 944
rect 35780 938 35786 944
rect 32400 820 32580 821
rect 36400 821 36401 999
rect 36579 821 36580 999
rect 39734 996 39740 1002
rect 39780 996 39786 1002
rect 39728 990 39734 996
rect 39786 990 39792 996
rect 39728 944 39734 950
rect 39786 944 39792 950
rect 39734 938 39740 944
rect 39780 938 39786 944
rect 36400 820 36580 821
rect 3262 808 3268 814
rect 3308 808 3314 814
rect 7262 808 7268 814
rect 7308 808 7314 814
rect 11262 808 11268 814
rect 11308 808 11314 814
rect 15262 808 15268 814
rect 15308 808 15314 814
rect 19262 808 19268 814
rect 19308 808 19314 814
rect 23262 808 23268 814
rect 23308 808 23314 814
rect 27262 808 27268 814
rect 27308 808 27314 814
rect 31262 808 31268 814
rect 31308 808 31314 814
rect 35262 808 35268 814
rect 35308 808 35314 814
rect 39262 808 39268 814
rect 39308 808 39314 814
rect 3256 802 3262 808
rect 3314 802 3320 808
rect 7256 802 7262 808
rect 7314 802 7320 808
rect 11256 802 11262 808
rect 11314 802 11320 808
rect 15256 802 15262 808
rect 15314 802 15320 808
rect 19256 802 19262 808
rect 19314 802 19320 808
rect 23256 802 23262 808
rect 23314 802 23320 808
rect 27256 802 27262 808
rect 27314 802 27320 808
rect 31256 802 31262 808
rect 31314 802 31320 808
rect 35256 802 35262 808
rect 35314 802 35320 808
rect 39256 802 39262 808
rect 39314 802 39320 808
rect 3256 756 3262 762
rect 3314 756 3320 762
rect 7256 756 7262 762
rect 7314 756 7320 762
rect 11256 756 11262 762
rect 11314 756 11320 762
rect 15256 756 15262 762
rect 15314 756 15320 762
rect 19256 756 19262 762
rect 19314 756 19320 762
rect 23256 756 23262 762
rect 23314 756 23320 762
rect 27256 756 27262 762
rect 27314 756 27320 762
rect 31256 756 31262 762
rect 31314 756 31320 762
rect 35256 756 35262 762
rect 35314 756 35320 762
rect 39256 756 39262 762
rect 39314 756 39320 762
rect 3262 750 3268 756
rect 3308 750 3314 756
rect 7262 750 7268 756
rect 7308 750 7314 756
rect 11262 750 11268 756
rect 11308 750 11314 756
rect 15262 750 15268 756
rect 15308 750 15314 756
rect 19262 750 19268 756
rect 19308 750 19314 756
rect 23262 750 23268 756
rect 23308 750 23314 756
rect 27262 750 27268 756
rect 27308 750 27314 756
rect 31262 750 31268 756
rect 31308 750 31314 756
rect 35262 750 35268 756
rect 35308 750 35314 756
rect 39262 750 39268 756
rect 39308 750 39314 756
rect 2240 296 2480 320
rect 2240 104 2264 296
rect 2456 104 2480 296
rect 2240 80 2480 104
rect 6240 296 6480 320
rect 6240 104 6264 296
rect 6456 104 6480 296
rect 6240 80 6480 104
rect 10240 296 10480 320
rect 10240 104 10264 296
rect 10456 104 10480 296
rect 10240 80 10480 104
rect 14240 296 14480 320
rect 14240 104 14264 296
rect 14456 104 14480 296
rect 14240 80 14480 104
rect 18240 296 18480 320
rect 18240 104 18264 296
rect 18456 104 18480 296
rect 18240 80 18480 104
rect 22240 296 22480 320
rect 22240 104 22264 296
rect 22456 104 22480 296
rect 22240 80 22480 104
rect 26240 296 26480 320
rect 26240 104 26264 296
rect 26456 104 26480 296
rect 26240 80 26480 104
rect 30240 296 30480 320
rect 30240 104 30264 296
rect 30456 104 30480 296
rect 30240 80 30480 104
rect 34240 296 34480 320
rect 34240 104 34264 296
rect 34456 104 34480 296
rect 34240 80 34480 104
rect 38240 296 38480 320
rect 38240 104 38264 296
rect 38456 104 38480 296
rect 38240 80 38480 104
use fgcell_amp_MiM_cap_1_5  fgcell_amp_MiM_cap_1_5_0
array 0 9 4000 0 9 3000
timestamp 1717597427
transform 1 0 -524 0 1 4198
box 458 -4198 4490 -1570
<< end >>
