magic
tech sky130A
magscale 1 2
timestamp 1716993393
<< error_p >>
rect 543 -2227 590 -1594
rect 597 -2281 644 -1648
rect 1234 -2292 1281 -1659
rect 1913 -1713 2008 -1694
rect 1288 -2346 1335 -1713
rect 1827 -1760 2008 -1713
rect 1913 -1818 2124 -1760
rect 1913 -2357 2037 -1818
rect 2113 -2191 2124 -1991
rect 1913 -2393 2026 -2357
rect 1979 -2411 2026 -2393
rect 2646 -2422 2663 -1806
rect 2700 -2471 2717 -1855
rect 3367 -2517 3384 -1901
rect 3421 -2566 3438 -1950
rect 4088 -2612 4105 -1996
rect 4142 -2661 4159 -2045
rect 4711 -2057 4826 -2045
rect 4718 -2091 4826 -2057
rect 4711 -2103 4826 -2091
rect 4768 -2158 4826 -2103
rect 4809 -2707 4826 -2158
rect 4827 -2158 4892 -2122
rect 4827 -2216 4978 -2158
rect 4827 -2707 4921 -2216
rect 4827 -2773 4892 -2707
rect 5500 -2802 5547 -2169
rect 5554 -2856 5601 -2223
rect 6191 -2867 6238 -2234
rect 6245 -2921 6292 -2288
use diffamp_nmos  x1
timestamp 1716993393
transform 1 0 65 0 1 2770
box -195 -5738 6900 200
<< end >>
