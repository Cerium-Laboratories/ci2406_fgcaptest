magic
tech sky130A
magscale 1 2
timestamp 1717598742
<< error_s >>
rect 64882 3800 65038 3960
rect 9770 -14600 9783 -14364
rect 20219 -14380 20243 -14364
rect 20243 -14600 20246 -14380
rect 24770 -14600 24783 -14364
rect 35219 -14380 35243 -14364
rect 35243 -14600 35246 -14380
rect 39770 -14520 39783 -14364
rect 50219 -14380 50243 -14364
rect 54770 -14380 54783 -14364
rect 65219 -14380 65243 -14364
rect 50243 -14600 50246 -14380
rect 54770 -14600 54783 -14520
rect 65243 -14600 65246 -14380
rect 69770 -14520 69783 -14364
rect 80219 -14380 80243 -14364
rect 80243 -14600 80246 -14380
rect 9451 -14688 9684 -14672
rect 24451 -14688 24684 -14672
rect 39451 -14688 39684 -14672
rect 54451 -14688 54684 -14672
rect 69451 -14688 69684 -14672
rect 9448 -14908 9451 -14688
rect 20551 -14742 20605 -14726
rect 20605 -14962 20608 -14742
rect 24448 -14908 24451 -14688
rect 35372 -14742 35605 -14726
rect 39448 -14742 39451 -14688
rect 50551 -14742 50605 -14726
rect 35605 -14962 35608 -14742
rect 50605 -14962 50608 -14742
rect 54448 -14908 54451 -14688
rect 65372 -14742 65605 -14726
rect 69448 -14742 69451 -14688
rect 80372 -14742 80605 -14726
rect 65605 -14962 65608 -14742
rect 80605 -14962 80608 -14742
rect 9141 -14998 9364 -14992
rect 24141 -14998 24364 -14992
rect 39141 -14998 39364 -14992
rect 54141 -14998 54364 -14992
rect 69141 -14998 69364 -14992
rect 9128 -15228 9141 -14998
rect 20861 -15056 20919 -15046
rect 20919 -15282 20928 -15056
rect 24128 -15228 24141 -14998
rect 35692 -15056 35919 -15046
rect 39128 -15056 39141 -14998
rect 50861 -15056 50919 -15046
rect 35919 -15282 35928 -15056
rect 50919 -15282 50928 -15056
rect 54128 -15228 54141 -14998
rect 65692 -15056 65919 -15046
rect 69128 -15056 69141 -14998
rect 80692 -15056 80919 -15046
rect 65919 -15282 65928 -15056
rect 80919 -15282 80928 -15056
rect 8811 -15328 9044 -15312
rect 23811 -15328 24044 -15312
rect 38811 -15328 39044 -15312
rect 53811 -15328 54044 -15312
rect 68811 -15328 69044 -15312
rect 8808 -15548 8811 -15328
rect 21191 -15382 21245 -15366
rect 21245 -15390 21248 -15382
rect 23808 -15390 23811 -15328
rect 36012 -15382 36245 -15366
rect 38808 -15382 38811 -15328
rect 51191 -15382 51245 -15366
rect 36245 -15390 36248 -15382
rect 51245 -15390 51248 -15382
rect 53808 -15390 53811 -15328
rect 66012 -15382 66245 -15366
rect 68808 -15382 68811 -15328
rect 81012 -15382 81245 -15366
rect 66245 -15390 66248 -15382
rect 81245 -15390 81248 -15382
rect 8497 -15642 8721 -15635
rect 23497 -15642 23721 -15635
rect 38497 -15642 38721 -15635
rect 53497 -15642 53721 -15635
rect 68497 -15642 68721 -15635
rect 8485 -15662 8497 -15642
rect 23485 -15662 23497 -15642
rect 38485 -15662 38497 -15642
rect 53485 -15662 53497 -15642
rect 68485 -15662 68497 -15642
rect 9943 -22517 9977 -22483
rect 9979 -22555 10015 -22483
rect 19985 -22555 20021 -22483
rect 20023 -22517 20057 -22483
rect 24943 -22517 24977 -22483
rect 24979 -22555 25015 -22483
rect 34985 -22555 35021 -22483
rect 35023 -22517 35057 -22483
rect 39943 -22517 39977 -22483
rect 39979 -22555 40015 -22483
rect 49985 -22555 50021 -22483
rect 50023 -22517 50057 -22483
rect 54943 -22517 54977 -22483
rect 54979 -22555 55015 -22483
rect 64985 -22555 65021 -22483
rect 65023 -22517 65057 -22483
rect 69943 -22517 69977 -22483
rect 69979 -22555 70015 -22483
rect 79985 -22555 80021 -22483
rect 80023 -22517 80057 -22483
rect 21514 -28109 21517 -28098
rect 36514 -28109 36517 -28098
rect 51514 -28109 51517 -28098
rect 66514 -28109 66517 -28098
rect 81514 -28109 81517 -28098
rect 21286 -28125 21514 -28109
rect 36286 -28125 36514 -28109
rect 51286 -28125 51514 -28109
rect 66286 -28125 66514 -28109
rect 81286 -28125 81514 -28109
rect 8754 -28378 8757 -28158
rect 23754 -28378 23757 -28158
rect 38754 -28378 38757 -28337
rect 53754 -28378 53757 -28158
rect 68754 -28378 68757 -28337
rect 8757 -28394 8990 -28378
rect 23757 -28380 23759 -28378
rect 38757 -28380 38759 -28378
rect 53757 -28380 53759 -28378
rect 68757 -28380 68759 -28378
rect 21191 -28432 21194 -28380
rect 23759 -28394 23990 -28380
rect 36191 -28432 36194 -28380
rect 38759 -28394 38811 -28380
rect 51191 -28432 51194 -28380
rect 53759 -28394 53990 -28380
rect 66191 -28432 66194 -28380
rect 68759 -28394 68811 -28380
rect 81191 -28432 81194 -28380
rect 20958 -28448 21191 -28432
rect 35958 -28448 36191 -28432
rect 50958 -28448 51191 -28432
rect 65958 -28448 66191 -28432
rect 80958 -28448 81191 -28432
rect 9074 -28698 9077 -28478
rect 24074 -28698 24077 -28478
rect 9077 -28714 9310 -28698
rect 20871 -28752 20874 -28698
rect 24077 -28714 24310 -28698
rect 35871 -28752 35874 -28532
rect 39074 -28698 39077 -28478
rect 54074 -28698 54077 -28478
rect 39077 -28714 39131 -28698
rect 50871 -28752 50874 -28698
rect 54077 -28714 54310 -28698
rect 65871 -28752 65874 -28532
rect 69074 -28698 69077 -28478
rect 69077 -28714 69131 -28698
rect 80871 -28752 80874 -28532
rect 20754 -28768 20871 -28752
rect 35754 -28768 35871 -28752
rect 50754 -28768 50871 -28752
rect 65754 -28768 65871 -28752
rect 80754 -28768 80871 -28752
rect 9394 -29018 9397 -28798
rect 24394 -29018 24397 -28798
rect 9397 -29034 9630 -29018
rect 20551 -29072 20554 -29018
rect 24397 -29034 24630 -29018
rect 35551 -29072 35554 -28869
rect 39394 -29018 39397 -28869
rect 54394 -29018 54397 -28798
rect 39397 -29034 39451 -29018
rect 50551 -29072 50554 -29018
rect 54397 -29034 54630 -29018
rect 65551 -29072 65554 -28869
rect 69394 -29018 69397 -28869
rect 69397 -29034 69451 -29018
rect 80551 -29072 80554 -28869
rect 20318 -29088 20551 -29072
rect 35318 -29088 35551 -29072
rect 50318 -29088 50551 -29072
rect 65318 -29088 65551 -29072
rect 80318 -29088 80551 -29072
rect 9756 -29380 9759 -29160
rect 24756 -29380 24759 -29160
rect 9759 -29396 9783 -29380
rect 20219 -29396 20232 -29380
rect 24759 -29396 24783 -29380
rect 35219 -29396 35232 -29160
rect 39756 -29380 39759 -29160
rect 54756 -29380 54759 -29160
rect 39759 -29396 39783 -29380
rect 50219 -29396 50232 -29380
rect 54759 -29396 54783 -29380
rect 65219 -29396 65232 -29160
rect 69756 -29380 69759 -29160
rect 69759 -29396 69783 -29380
rect 80219 -29396 80232 -29160
<< metal1 >>
rect 64882 3960 65038 3966
rect 51996 3954 64882 3960
rect 51996 3902 52028 3954
rect 52132 3902 53628 3954
rect 53732 3902 55228 3954
rect 55332 3902 56828 3954
rect 56932 3902 58428 3954
rect 58532 3902 60028 3954
rect 60132 3902 61628 3954
rect 61732 3902 63228 3954
rect 63332 3902 64882 3954
rect 51996 3800 64882 3902
rect 52360 3708 52476 3714
rect 52360 3604 52366 3708
rect 52470 3604 52476 3708
rect 52746 3688 52830 3800
rect 53160 3708 53276 3714
rect 52360 3598 52476 3604
rect 53160 3604 53166 3708
rect 53270 3604 53276 3708
rect 53546 3688 53630 3800
rect 53960 3708 54076 3714
rect 53160 3598 53276 3604
rect 53960 3604 53966 3708
rect 54070 3604 54076 3708
rect 54346 3688 54430 3800
rect 54760 3708 54876 3714
rect 53960 3598 54076 3604
rect 54760 3604 54766 3708
rect 54870 3604 54876 3708
rect 55146 3688 55230 3800
rect 55560 3708 55676 3714
rect 54760 3598 54876 3604
rect 55560 3604 55566 3708
rect 55670 3604 55676 3708
rect 55946 3688 56030 3800
rect 56360 3708 56476 3714
rect 55560 3598 55676 3604
rect 56360 3604 56366 3708
rect 56470 3604 56476 3708
rect 56746 3688 56830 3800
rect 57160 3708 57276 3714
rect 56360 3598 56476 3604
rect 57160 3604 57166 3708
rect 57270 3604 57276 3708
rect 57546 3688 57630 3800
rect 57960 3708 58076 3714
rect 57160 3598 57276 3604
rect 57960 3604 57966 3708
rect 58070 3604 58076 3708
rect 58346 3688 58430 3800
rect 58760 3708 58876 3714
rect 57960 3598 58076 3604
rect 58760 3604 58766 3708
rect 58870 3604 58876 3708
rect 59146 3688 59230 3800
rect 59560 3708 59676 3714
rect 58760 3598 58876 3604
rect 59560 3604 59566 3708
rect 59670 3604 59676 3708
rect 59946 3688 60030 3800
rect 60360 3708 60476 3714
rect 59560 3598 59676 3604
rect 60360 3604 60366 3708
rect 60470 3604 60476 3708
rect 60746 3688 60830 3800
rect 61160 3708 61276 3714
rect 60360 3598 60476 3604
rect 61160 3604 61166 3708
rect 61270 3604 61276 3708
rect 61546 3688 61630 3800
rect 61960 3708 62076 3714
rect 61160 3598 61276 3604
rect 61960 3604 61966 3708
rect 62070 3604 62076 3708
rect 62346 3688 62430 3800
rect 62760 3708 62876 3714
rect 61960 3598 62076 3604
rect 62760 3604 62766 3708
rect 62870 3604 62876 3708
rect 63146 3688 63230 3800
rect 63560 3708 63676 3714
rect 62760 3598 62876 3604
rect 63560 3604 63566 3708
rect 63670 3604 63676 3708
rect 63946 3688 64030 3800
rect 64360 3708 64476 3714
rect 63560 3598 63676 3604
rect 64360 3604 64366 3708
rect 64470 3604 64476 3708
rect 64746 3688 64830 3800
rect 64882 3794 65038 3800
rect 64360 3598 64476 3604
rect 106000 -20440 106260 -20400
rect 106000 -27780 106020 -20440
rect 106220 -27780 106260 -20440
rect 106000 -27820 106260 -27780
<< via1 >>
rect 52028 4260 52132 4312
rect 53628 4260 53732 4312
rect 55228 4260 55332 4312
rect 56828 4260 56932 4312
rect 58428 4260 58532 4312
rect 60028 4260 60132 4312
rect 61628 4260 61732 4312
rect 63228 4260 63332 4312
rect 52028 3902 52132 3954
rect 53628 3902 53732 3954
rect 55228 3902 55332 3954
rect 56828 3902 56932 3954
rect 58428 3902 58532 3954
rect 60028 3902 60132 3954
rect 61628 3902 61732 3954
rect 63228 3902 63332 3954
rect 64882 3800 65038 3960
rect 52366 3604 52470 3708
rect 53166 3604 53270 3708
rect 53966 3604 54070 3708
rect 54766 3604 54870 3708
rect 55566 3604 55670 3708
rect 56366 3604 56470 3708
rect 57166 3604 57270 3708
rect 57966 3604 58070 3708
rect 58766 3604 58870 3708
rect 59566 3604 59670 3708
rect 60366 3604 60470 3708
rect 61166 3604 61270 3708
rect 61966 3604 62070 3708
rect 62766 3604 62870 3708
rect 63566 3604 63670 3708
rect 64366 3604 64470 3708
rect 106020 -27780 106220 -20440
<< metal2 >>
rect 52022 4312 52138 4318
rect 52022 4260 52028 4312
rect 52132 4260 52138 4312
rect 52022 3954 52138 4260
rect 53622 4312 53738 4318
rect 53622 4260 53628 4312
rect 53732 4260 53738 4312
rect 52022 3902 52028 3954
rect 52132 3902 52138 3954
rect 52022 3896 52138 3902
rect 52360 3708 52476 4000
rect 52360 3604 52366 3708
rect 52470 3604 52476 3708
rect 52360 3598 52476 3604
rect 53160 3708 53276 4000
rect 53622 3954 53738 4260
rect 55222 4312 55338 4318
rect 55222 4260 55228 4312
rect 55332 4260 55338 4312
rect 53622 3902 53628 3954
rect 53732 3902 53738 3954
rect 53622 3896 53738 3902
rect 53160 3604 53166 3708
rect 53270 3604 53276 3708
rect 53160 3598 53276 3604
rect 53960 3708 54076 4000
rect 53960 3604 53966 3708
rect 54070 3604 54076 3708
rect 53960 3598 54076 3604
rect 54760 3708 54876 4000
rect 55222 3954 55338 4260
rect 56822 4312 56938 4318
rect 56822 4260 56828 4312
rect 56932 4260 56938 4312
rect 55222 3902 55228 3954
rect 55332 3902 55338 3954
rect 55222 3896 55338 3902
rect 54760 3604 54766 3708
rect 54870 3604 54876 3708
rect 54760 3598 54876 3604
rect 55560 3708 55676 4000
rect 55560 3604 55566 3708
rect 55670 3604 55676 3708
rect 55560 3598 55676 3604
rect 56360 3708 56476 4000
rect 56822 3954 56938 4260
rect 58422 4312 58538 4318
rect 58422 4260 58428 4312
rect 58532 4260 58538 4312
rect 56822 3902 56828 3954
rect 56932 3902 56938 3954
rect 56822 3896 56938 3902
rect 56360 3604 56366 3708
rect 56470 3604 56476 3708
rect 56360 3598 56476 3604
rect 57160 3708 57276 4000
rect 57160 3604 57166 3708
rect 57270 3604 57276 3708
rect 57160 3598 57276 3604
rect 57960 3708 58076 4000
rect 58422 3954 58538 4260
rect 60022 4312 60138 4318
rect 60022 4260 60028 4312
rect 60132 4260 60138 4312
rect 58422 3902 58428 3954
rect 58532 3902 58538 3954
rect 58422 3896 58538 3902
rect 57960 3604 57966 3708
rect 58070 3604 58076 3708
rect 57960 3598 58076 3604
rect 58760 3708 58876 4000
rect 58760 3604 58766 3708
rect 58870 3604 58876 3708
rect 58760 3598 58876 3604
rect 59560 3708 59676 4000
rect 60022 3954 60138 4260
rect 61622 4312 61738 4318
rect 61622 4260 61628 4312
rect 61732 4260 61738 4312
rect 60022 3902 60028 3954
rect 60132 3902 60138 3954
rect 60022 3896 60138 3902
rect 59560 3604 59566 3708
rect 59670 3604 59676 3708
rect 59560 3598 59676 3604
rect 60360 3708 60476 4000
rect 60360 3604 60366 3708
rect 60470 3604 60476 3708
rect 60360 3598 60476 3604
rect 61160 3708 61276 4000
rect 61622 3954 61738 4260
rect 63222 4312 63338 4318
rect 63222 4260 63228 4312
rect 63332 4260 63338 4312
rect 61622 3902 61628 3954
rect 61732 3902 61738 3954
rect 61622 3896 61738 3902
rect 61160 3604 61166 3708
rect 61270 3604 61276 3708
rect 61160 3598 61276 3604
rect 61960 3708 62076 4000
rect 61960 3604 61966 3708
rect 62070 3604 62076 3708
rect 61960 3598 62076 3604
rect 62760 3708 62876 4000
rect 63222 3954 63338 4260
rect 63222 3902 63228 3954
rect 63332 3902 63338 3954
rect 63222 3896 63338 3902
rect 62760 3604 62766 3708
rect 62870 3604 62876 3708
rect 62760 3598 62876 3604
rect 63560 3708 63676 4000
rect 63560 3604 63566 3708
rect 63670 3604 63676 3708
rect 63560 3598 63676 3604
rect 64360 3708 64476 4000
rect 64882 3960 65038 4260
rect 64882 3794 65038 3800
rect 64360 3604 64366 3708
rect 64470 3604 64476 3708
rect 64360 3598 64476 3604
rect 106000 -20440 106260 -20400
rect 106000 -27780 106020 -20440
rect 106220 -27780 106260 -20440
rect 106000 -27820 106260 -27780
<< via2 >>
rect 106020 -27780 106220 -20440
<< metal3 >>
rect 48200 91000 49800 91200
rect 52200 91000 53800 91200
rect 54600 91000 55000 91200
rect 55800 91000 56200 91200
rect 57000 91000 57400 91200
rect 58200 91000 58600 91200
rect 59400 91000 59800 91200
rect 60600 91000 61000 91200
rect 61800 91000 62200 91200
rect 63000 91000 63400 91200
rect 64200 91000 64600 91200
rect 65400 91000 67000 91200
rect 69400 91000 71000 91200
rect 14400 -4820 45500 -4800
rect 14400 -5980 14420 -4820
rect 15580 -5980 45500 -4820
rect 14400 -6000 45500 -5980
rect 45720 -6200 47040 -5200
rect 29400 -6220 47040 -6200
rect 29400 -7380 29420 -6220
rect 30580 -7380 47040 -6220
rect 29400 -7400 47040 -7380
rect 48800 -7800 49600 -5200
rect 44400 -7820 49600 -7800
rect 44400 -8580 44420 -7820
rect 45580 -8580 49600 -7820
rect 44400 -8600 49600 -8580
rect 74400 -7820 75600 -5200
rect 87800 -5240 92200 -5200
rect 87800 -5760 87840 -5240
rect 92160 -5760 92200 -5240
rect 87800 -5800 92200 -5760
rect 74400 -8580 74420 -7820
rect 75580 -8580 75600 -7820
rect 74400 -8620 75600 -8580
rect 95920 -20440 106260 -20400
rect 95920 -27780 106020 -20440
rect 106220 -27780 106260 -20440
rect 95920 -27820 106260 -27780
<< via3 >>
rect 14420 -5980 15580 -4820
rect 29420 -7380 30580 -6220
rect 44420 -8580 45580 -7820
rect 87840 -5760 92160 -5240
rect 74420 -8580 75580 -7820
<< metal4 >>
rect 14400 -4820 15600 -4800
rect 14400 -5980 14420 -4820
rect 15580 -5980 15600 -4820
rect 14400 -8810 15600 -5980
rect 29400 -6220 30600 -6200
rect 29400 -7380 29420 -6220
rect 30580 -7380 30600 -6220
rect 29400 -8810 30600 -7380
rect 44400 -7820 45600 -7800
rect 44400 -8580 44420 -7820
rect 45580 -8580 45600 -7820
rect 44400 -8820 45600 -8580
rect 58000 -9000 62000 -5200
rect 87800 -5240 92200 -5200
rect 87800 -5760 87840 -5240
rect 92160 -5760 92200 -5240
rect 87800 -5800 92200 -5760
rect 74400 -7820 75600 -7800
rect 74400 -8580 74420 -7820
rect 75580 -8580 75600 -7820
rect 74400 -8820 75600 -8580
rect 58160 -13800 61878 -9000
<< via4 >>
rect 87840 -5760 92160 -5240
<< metal5 >>
rect -1000 -29957 -200 -3000
rect 87800 -5240 92200 -5200
rect 87800 -5760 87840 -5240
rect 92160 -5760 92200 -5240
rect 87800 -14600 92200 -5760
rect 108800 -14020 113200 -5200
rect 9510 -28396 20500 -15374
rect 24510 -28396 35500 -15374
rect 39510 -28396 50500 -15374
rect 54510 -28396 65500 -15374
rect 69510 -28396 80500 -15374
rect 83720 -29160 96280 -14600
rect 104720 -29160 117280 -14600
rect -1000 -34800 7500 -29957
rect 83460 -29960 96540 -29420
rect 82500 -30800 96540 -29960
rect 120120 -30800 120920 -2000
rect 82500 -34800 120920 -30800
use array_core  array_core_0
timestamp 1717598570
transform 1 0 40000 0 1 0
box -41000 -5200 80920 91200
use bare_pad_gnd  bare_pad_gnd_0
timestamp 1717393140
transform 1 0 83460 0 1 -29420
box 0 0 13080 15080
use pad_minesd_short  pad_minesd_short_0
timestamp 1717582298
transform -1 0 37500 0 -1 5200
box 0 14007 15000 40000
use pad_minesd_short  pad_minesd_short_1
timestamp 1717582298
transform -1 0 22500 0 -1 5200
box 0 14007 15000 40000
use pad_minesd_short  pad_minesd_short_2
timestamp 1717582298
transform -1 0 67500 0 -1 5200
box 0 14007 15000 40000
use pad_minesd_short  pad_minesd_short_3
timestamp 1717582298
transform -1 0 52500 0 -1 5200
box 0 14007 15000 40000
use pad_minesd_short  pad_minesd_short_4
timestamp 1717582298
transform -1 0 82500 0 -1 5200
box 0 14007 15000 40000
use vtun_pad  vtun_pad_0
timestamp 1717596487
transform 1 0 104460 0 1 -29420
box 0 0 13080 16200
<< labels >>
flabel metal5 83720 -29160 96280 -14600 0 FreeSans 6400 0 0 0 VGND
flabel metal5 39510 -28396 50500 -15374 0 FreeSans 6400 0 0 0 VOUT0
flabel metal5 69510 -28396 80500 -15374 0 FreeSans 6400 0 0 0 VOUT1
flabel metal5 54510 -28396 65500 -15374 0 FreeSans 6400 0 0 0 VINJ
flabel metal5 24510 -28396 35500 -15374 0 FreeSans 6400 0 0 0 VCTRL
flabel metal5 9510 -28396 20500 -15374 0 FreeSans 6400 0 0 0 VSRC
flabel metal5 104720 -29160 117280 -14600 0 FreeSans 6400 0 0 0 VTUN
flabel metal3 54600 91000 55000 91200 0 FreeSans 800 0 0 0 addr[0]
port 3 n signal input
flabel metal3 55800 91000 56200 91200 0 FreeSans 800 0 0 0 addr[1]
port 4 n signal input
flabel metal3 57000 91000 57400 91200 0 FreeSans 800 0 0 0 addr[2]
port 5 n signal input
flabel metal3 58200 91000 58600 91200 0 FreeSans 800 0 0 0 addr[3]
port 6 n signal input
flabel metal3 59400 91000 59800 91200 0 FreeSans 800 0 0 0 addr[4]
port 7 n signal input
flabel metal3 60600 91000 61000 91200 0 FreeSans 800 0 0 0 addr[5]
port 8 n signal input
flabel metal3 61800 91000 62200 91200 0 FreeSans 800 0 0 0 addr[6]
port 9 n signal input
flabel metal3 63000 91000 63400 91200 0 FreeSans 800 0 0 0 addr[7]
port 10 n signal input
flabel metal3 64200 91000 64600 91200 0 FreeSans 800 0 0 0 addr[8]
port 11 n signal input
flabel metal3 52200 91000 53800 91200 0 FreeSans 1600 0 0 0 vssd2
port 2 n ground default
flabel metal3 65400 91000 67000 91200 0 FreeSans 1600 0 0 0 vccd2
port 1 n power default
flabel metal3 48200 91000 49800 91200 0 FreeSans 1600 0 0 0 vccd2
port 1 n power default
flabel metal3 69400 91000 71000 91200 0 FreeSans 1600 0 0 0 vssd2
port 2 n ground default
<< properties >>
string FIXED_BBOX -2000 -35800 121920 92200
<< end >>
