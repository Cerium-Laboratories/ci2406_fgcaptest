magic
tech sky130A
timestamp 1717034485
<< end >>
