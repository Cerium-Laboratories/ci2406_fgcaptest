magic
tech sky130A
magscale 1 2
timestamp 1717562480
<< pwell >>
rect -4843 -3702 4843 3702
<< psubdiff >>
rect -4807 3632 -4711 3666
rect 4711 3632 4807 3666
rect -4807 3570 -4773 3632
rect 4773 3570 4807 3632
rect -4807 -3632 -4773 -3570
rect 4773 -3632 4807 -3570
rect -4807 -3666 -4711 -3632
rect 4711 -3666 4807 -3632
<< psubdiffcont >>
rect -4711 3632 4711 3666
rect -4807 -3570 -4773 3570
rect 4773 -3570 4807 3570
rect -4711 -3666 4711 -3632
<< xpolycontact >>
rect 4395 3104 4677 3536
rect -4677 -3536 -4395 -3104
<< xpolyres >>
rect -4677 2718 -4017 3000
rect -4677 -3104 -4395 2718
rect -4299 -2718 -4017 2718
rect -3921 2718 -3261 3000
rect -3921 -2718 -3639 2718
rect -4299 -3000 -3639 -2718
rect -3543 -2718 -3261 2718
rect -3165 2718 -2505 3000
rect -3165 -2718 -2883 2718
rect -3543 -3000 -2883 -2718
rect -2787 -2718 -2505 2718
rect -2409 2718 -1749 3000
rect -2409 -2718 -2127 2718
rect -2787 -3000 -2127 -2718
rect -2031 -2718 -1749 2718
rect -1653 2718 -993 3000
rect -1653 -2718 -1371 2718
rect -2031 -3000 -1371 -2718
rect -1275 -2718 -993 2718
rect -897 2718 -237 3000
rect -897 -2718 -615 2718
rect -1275 -3000 -615 -2718
rect -519 -2718 -237 2718
rect -141 2718 519 3000
rect -141 -2718 141 2718
rect -519 -3000 141 -2718
rect 237 -2718 519 2718
rect 615 2718 1275 3000
rect 615 -2718 897 2718
rect 237 -3000 897 -2718
rect 993 -2718 1275 2718
rect 1371 2718 2031 3000
rect 1371 -2718 1653 2718
rect 993 -3000 1653 -2718
rect 1749 -2718 2031 2718
rect 2127 2718 2787 3000
rect 2127 -2718 2409 2718
rect 1749 -3000 2409 -2718
rect 2505 -2718 2787 2718
rect 2883 2718 3543 3000
rect 2883 -2718 3165 2718
rect 2505 -3000 3165 -2718
rect 3261 -2718 3543 2718
rect 3639 2718 4299 3000
rect 3639 -2718 3921 2718
rect 3261 -3000 3921 -2718
rect 4017 -2718 4299 2718
rect 4395 -2718 4677 3104
rect 4017 -3000 4677 -2718
<< locali >>
rect -4807 3632 -4711 3666
rect 4711 3632 4807 3666
rect -4807 3570 -4773 3632
rect 4773 3570 4807 3632
rect -4807 -3632 -4773 -3570
rect 4773 -3632 4807 -3570
rect -4807 -3666 -4711 -3632
rect 4711 -3666 4807 -3632
<< properties >>
string FIXED_BBOX -4790 -3649 4790 3649
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 30.0 m 1 nx 25 wmin 1.410 lmin 0.50 rho 2000 val 1.112meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
