magic
tech sky130A
magscale 1 2
timestamp 1717630197
<< pwell >>
rect 1700 1440 11386 9104
<< psubdiff >>
rect 1736 9034 1832 9068
rect 11254 9034 11350 9068
rect 1736 8972 1770 9034
rect 11316 8972 11350 9034
rect 1736 1510 1770 1572
rect 11316 1510 11350 1572
rect 1736 1476 1832 1510
rect 11254 1476 11350 1510
<< psubdiffcont >>
rect 1832 9034 11254 9068
rect 1736 1572 1770 8972
rect 11316 1572 11350 8972
rect 1832 1476 11254 1510
<< poly >>
rect 5600 10984 6030 11000
rect 5600 9616 5616 10984
rect 5650 9616 6030 10984
rect 5600 9600 6030 9616
rect 10830 10984 11260 11000
rect 10830 9616 11210 10984
rect 11244 9616 11260 10984
rect 10830 9600 11260 9616
<< polycont >>
rect 5616 9616 5650 10984
rect 11210 9616 11244 10984
<< xpolycontact >>
rect 10938 8406 11220 8938
rect 1866 1606 2148 2198
<< npolyres >>
rect 6030 9600 10830 11000
<< xpolyres >>
rect 1866 8020 2526 8302
rect 1866 2198 2148 8020
rect 2244 2584 2526 8020
rect 2622 8020 3282 8302
rect 2622 2584 2904 8020
rect 2244 2302 2904 2584
rect 3000 2584 3282 8020
rect 3378 8020 4038 8302
rect 3378 2584 3660 8020
rect 3000 2302 3660 2584
rect 3756 2584 4038 8020
rect 4134 8020 4794 8302
rect 4134 2584 4416 8020
rect 3756 2302 4416 2584
rect 4512 2584 4794 8020
rect 4890 8020 5550 8302
rect 4890 2584 5172 8020
rect 4512 2302 5172 2584
rect 5268 2584 5550 8020
rect 5646 8020 6306 8302
rect 5646 2584 5928 8020
rect 5268 2302 5928 2584
rect 6024 2584 6306 8020
rect 6402 8020 7062 8302
rect 6402 2584 6684 8020
rect 6024 2302 6684 2584
rect 6780 2584 7062 8020
rect 7158 8020 7818 8302
rect 7158 2584 7440 8020
rect 6780 2302 7440 2584
rect 7536 2584 7818 8020
rect 7914 8020 8574 8302
rect 7914 2584 8196 8020
rect 7536 2302 8196 2584
rect 8292 2584 8574 8020
rect 8670 8020 9330 8302
rect 8670 2584 8952 8020
rect 8292 2302 8952 2584
rect 9048 2584 9330 8020
rect 9426 8020 10086 8302
rect 9426 2584 9708 8020
rect 9048 2302 9708 2584
rect 9804 2584 10086 8020
rect 10182 8020 10842 8302
rect 10182 2584 10464 8020
rect 9804 2302 10464 2584
rect 10560 2584 10842 8020
rect 10938 2584 11220 8406
rect 10560 2302 11220 2584
<< locali >>
rect 5616 10984 5650 11000
rect 11210 10984 11244 11000
rect 5616 9600 5650 9616
rect 11210 9600 11244 9616
rect 1736 9034 1832 9068
rect 11254 9034 11350 9068
rect 1736 8972 1770 9034
rect 11316 8972 11350 9034
rect 1736 1510 1770 1572
rect 11316 1510 11350 1572
rect 1736 1476 1832 1510
rect 11254 1476 11350 1510
<< viali >>
rect 5616 9616 5650 10984
rect 5650 9616 6013 10984
rect 10847 9616 11210 10984
rect 11210 9616 11244 10984
rect 10920 8938 11220 8940
rect 10920 8406 10938 8938
rect 10938 8406 11220 8938
rect 10920 8400 11220 8406
rect 1866 1606 2148 2198
<< metal1 >>
rect 10800 11200 13080 11220
rect 4400 10984 6020 11000
rect 4400 10980 5616 10984
rect 4400 9620 4420 10980
rect 4400 9616 5616 9620
rect 6013 9616 6020 10984
rect 4400 9600 6020 9616
rect 10800 10984 12820 11200
rect 10800 9616 10847 10984
rect 11244 9616 12820 10984
rect 1700 9000 9800 9104
rect 1700 2220 1800 9000
rect 10800 8940 12820 9616
rect 10800 8400 10920 8940
rect 11220 8400 12820 8940
rect 10800 8200 12820 8400
rect 13060 8200 13080 11200
rect 10800 8180 13080 8200
rect 1700 2198 2160 2220
rect 1700 1606 1866 2198
rect 2148 1606 2160 2198
rect 1700 1540 2160 1606
rect 11280 1540 11380 7680
rect 1700 1440 11380 1540
<< via1 >>
rect 4420 9620 5616 10980
rect 5616 9620 6000 10980
rect 12820 8200 13060 11200
<< metal2 >>
rect 12800 11200 13080 11220
rect 4400 10980 6020 11000
rect 4400 9620 4420 10980
rect 6000 9620 6020 10980
rect 4400 9600 6020 9620
rect 12800 8200 12820 11200
rect 13060 8200 13080 11200
rect 12800 8180 13080 8200
<< via2 >>
rect 4420 9620 6000 10980
rect 12820 8200 13060 11200
<< metal3 >>
rect 4400 16160 8600 16200
rect 4400 15440 4440 16160
rect 8560 15440 8600 16160
rect 4400 15400 8600 15440
rect 4400 10980 6200 15400
rect 4400 9620 4420 10980
rect 6000 9620 6200 10980
rect 4400 9600 6200 9620
rect 12800 11200 13080 11220
rect 12800 8200 12820 11200
rect 13060 8200 13080 11200
rect 12800 8180 13080 8200
<< via3 >>
rect 4440 15440 8560 16160
rect 12820 8200 13060 11200
<< metal4 >>
rect 4400 16160 8600 16200
rect 4400 15440 4440 16160
rect 8560 15440 8600 16160
rect 4400 15400 8600 15440
rect 0 15056 13080 15080
rect 0 14820 24 15056
rect 260 14820 502 15056
rect 738 14820 822 15056
rect 1058 14820 1142 15056
rect 1378 14820 1462 15056
rect 1698 14820 1782 15056
rect 2018 14820 2102 15056
rect 2338 14820 2422 15056
rect 2658 14820 2742 15056
rect 2978 14820 3062 15056
rect 3298 14820 3382 15056
rect 3618 14820 3702 15056
rect 3938 14820 4022 15056
rect 4258 14820 4342 15056
rect 4578 14820 4662 15056
rect 4898 14820 4982 15056
rect 5218 14820 5302 15056
rect 5538 14820 5622 15056
rect 5858 14820 5942 15056
rect 6178 14820 6262 15056
rect 6498 14820 6582 15056
rect 6818 14820 6902 15056
rect 7138 14820 7222 15056
rect 7458 14820 7542 15056
rect 7778 14820 7862 15056
rect 8098 14820 8182 15056
rect 8418 14820 8502 15056
rect 8738 14820 8822 15056
rect 9058 14820 9142 15056
rect 9378 14820 9462 15056
rect 9698 14820 9782 15056
rect 10018 14820 10102 15056
rect 10338 14820 10422 15056
rect 10658 14820 10742 15056
rect 10978 14820 11062 15056
rect 11298 14820 11382 15056
rect 11618 14820 11702 15056
rect 11938 14820 12022 15056
rect 12258 14820 12342 15056
rect 12578 14820 12820 15056
rect 13056 14820 13080 15056
rect 0 14698 13080 14820
rect 0 14462 24 14698
rect 260 14462 12820 14698
rect 13056 14462 13080 14698
rect 0 14378 13080 14462
rect 0 14142 24 14378
rect 260 14142 12820 14378
rect 13056 14142 13080 14378
rect 0 14058 13080 14142
rect 0 13822 24 14058
rect 260 13822 12820 14058
rect 13056 13822 13080 14058
rect 0 13738 13080 13822
rect 0 13502 24 13738
rect 260 13502 12820 13738
rect 13056 13502 13080 13738
rect 0 13418 13080 13502
rect 0 13182 24 13418
rect 260 13182 12820 13418
rect 13056 13182 13080 13418
rect 0 13098 13080 13182
rect 0 12862 24 13098
rect 260 12862 12820 13098
rect 13056 12862 13080 13098
rect 0 12778 13080 12862
rect 0 12542 24 12778
rect 260 12542 12820 12778
rect 13056 12542 13080 12778
rect 0 12458 13080 12542
rect 0 12222 24 12458
rect 260 12222 12820 12458
rect 13056 12222 13080 12458
rect 0 12138 13080 12222
rect 0 11902 24 12138
rect 260 11902 12820 12138
rect 13056 11902 13080 12138
rect 0 11818 13080 11902
rect 0 11582 24 11818
rect 260 11582 12820 11818
rect 13056 11582 13080 11818
rect 0 11498 13080 11582
rect 0 11262 24 11498
rect 260 11262 12820 11498
rect 13056 11262 13080 11498
rect 0 11200 13080 11262
rect 0 11178 12820 11200
rect 0 10942 24 11178
rect 260 10942 12820 11178
rect 0 10858 12820 10942
rect 0 10622 24 10858
rect 260 10622 12820 10858
rect 0 10538 12820 10622
rect 0 10302 24 10538
rect 260 10302 12820 10538
rect 0 10218 12820 10302
rect 0 9982 24 10218
rect 260 9982 12820 10218
rect 0 9898 12820 9982
rect 0 9662 24 9898
rect 260 9662 12820 9898
rect 0 9578 12820 9662
rect 0 9342 24 9578
rect 260 9342 12820 9578
rect 0 9258 12820 9342
rect 0 9022 24 9258
rect 260 9022 12820 9258
rect 0 8938 12820 9022
rect 0 8702 24 8938
rect 260 8702 12820 8938
rect 0 8618 12820 8702
rect 0 8382 24 8618
rect 260 8382 12820 8618
rect 0 8298 12820 8382
rect 0 8062 24 8298
rect 260 8062 12820 8298
rect 13060 8200 13080 11200
rect 13056 8062 13080 8200
rect 0 7978 13080 8062
rect 0 7742 24 7978
rect 260 7742 12820 7978
rect 13056 7742 13080 7978
rect 0 7658 13080 7742
rect 0 7422 24 7658
rect 260 7422 12820 7658
rect 13056 7422 13080 7658
rect 0 7338 13080 7422
rect 0 7102 24 7338
rect 260 7102 12820 7338
rect 13056 7102 13080 7338
rect 0 7018 13080 7102
rect 0 6782 24 7018
rect 260 6782 12820 7018
rect 13056 6782 13080 7018
rect 0 6698 13080 6782
rect 0 6462 24 6698
rect 260 6462 12820 6698
rect 13056 6462 13080 6698
rect 0 6378 13080 6462
rect 0 6142 24 6378
rect 260 6142 12820 6378
rect 13056 6142 13080 6378
rect 0 6058 13080 6142
rect 0 5822 24 6058
rect 260 5822 12820 6058
rect 13056 5822 13080 6058
rect 0 5738 13080 5822
rect 0 5502 24 5738
rect 260 5502 12820 5738
rect 13056 5502 13080 5738
rect 0 5418 13080 5502
rect 0 5182 24 5418
rect 260 5182 12820 5418
rect 13056 5182 13080 5418
rect 0 5098 13080 5182
rect 0 4862 24 5098
rect 260 4862 12820 5098
rect 13056 4862 13080 5098
rect 0 4778 13080 4862
rect 0 4542 24 4778
rect 260 4542 12820 4778
rect 13056 4542 13080 4778
rect 0 4458 13080 4542
rect 0 4222 24 4458
rect 260 4222 12820 4458
rect 13056 4222 13080 4458
rect 0 4138 13080 4222
rect 0 3902 24 4138
rect 260 3902 12820 4138
rect 13056 3902 13080 4138
rect 0 3818 13080 3902
rect 0 3582 24 3818
rect 260 3582 12820 3818
rect 13056 3582 13080 3818
rect 0 3498 13080 3582
rect 0 3262 24 3498
rect 260 3262 12820 3498
rect 13056 3262 13080 3498
rect 0 3178 13080 3262
rect 0 2942 24 3178
rect 260 2942 12820 3178
rect 13056 2942 13080 3178
rect 0 2858 13080 2942
rect 0 2622 24 2858
rect 260 2622 12820 2858
rect 13056 2622 13080 2858
rect 0 2538 13080 2622
rect 0 2302 24 2538
rect 260 2302 12820 2538
rect 13056 2302 13080 2538
rect 0 2218 13080 2302
rect 0 1982 24 2218
rect 260 1982 12820 2218
rect 13056 1982 13080 2218
rect 0 1898 13080 1982
rect 0 1662 24 1898
rect 260 1662 12820 1898
rect 13056 1662 13080 1898
rect 0 1578 13080 1662
rect 0 1342 24 1578
rect 260 1342 12820 1578
rect 13056 1342 13080 1578
rect 0 1258 13080 1342
rect 0 1022 24 1258
rect 260 1022 12820 1258
rect 13056 1022 13080 1258
rect 0 938 13080 1022
rect 0 702 24 938
rect 260 702 12820 938
rect 13056 702 13080 938
rect 0 618 13080 702
rect 0 382 24 618
rect 260 382 12820 618
rect 13056 382 13080 618
rect 0 260 13080 382
rect 0 24 24 260
rect 260 24 502 260
rect 738 24 822 260
rect 1058 24 1142 260
rect 1378 24 1462 260
rect 1698 24 1782 260
rect 2018 24 2102 260
rect 2338 24 2422 260
rect 2658 24 2742 260
rect 2978 24 3062 260
rect 3298 24 3382 260
rect 3618 24 3702 260
rect 3938 24 4022 260
rect 4258 24 4342 260
rect 4578 24 4662 260
rect 4898 24 4982 260
rect 5218 24 5302 260
rect 5538 24 5622 260
rect 5858 24 5942 260
rect 6178 24 6262 260
rect 6498 24 6582 260
rect 6818 24 6902 260
rect 7138 24 7222 260
rect 7458 24 7542 260
rect 7778 24 7862 260
rect 8098 24 8182 260
rect 8418 24 8502 260
rect 8738 24 8822 260
rect 9058 24 9142 260
rect 9378 24 9462 260
rect 9698 24 9782 260
rect 10018 24 10102 260
rect 10338 24 10422 260
rect 10658 24 10742 260
rect 10978 24 11062 260
rect 11298 24 11382 260
rect 11618 24 11702 260
rect 11938 24 12022 260
rect 12258 24 12342 260
rect 12578 24 12820 260
rect 13056 24 13080 260
rect 0 0 13080 24
<< via4 >>
rect 24 14820 260 15056
rect 502 14820 738 15056
rect 822 14820 1058 15056
rect 1142 14820 1378 15056
rect 1462 14820 1698 15056
rect 1782 14820 2018 15056
rect 2102 14820 2338 15056
rect 2422 14820 2658 15056
rect 2742 14820 2978 15056
rect 3062 14820 3298 15056
rect 3382 14820 3618 15056
rect 3702 14820 3938 15056
rect 4022 14820 4258 15056
rect 4342 14820 4578 15056
rect 4662 14820 4898 15056
rect 4982 14820 5218 15056
rect 5302 14820 5538 15056
rect 5622 14820 5858 15056
rect 5942 14820 6178 15056
rect 6262 14820 6498 15056
rect 6582 14820 6818 15056
rect 6902 14820 7138 15056
rect 7222 14820 7458 15056
rect 7542 14820 7778 15056
rect 7862 14820 8098 15056
rect 8182 14820 8418 15056
rect 8502 14820 8738 15056
rect 8822 14820 9058 15056
rect 9142 14820 9378 15056
rect 9462 14820 9698 15056
rect 9782 14820 10018 15056
rect 10102 14820 10338 15056
rect 10422 14820 10658 15056
rect 10742 14820 10978 15056
rect 11062 14820 11298 15056
rect 11382 14820 11618 15056
rect 11702 14820 11938 15056
rect 12022 14820 12258 15056
rect 12342 14820 12578 15056
rect 12820 14820 13056 15056
rect 24 14462 260 14698
rect 12820 14462 13056 14698
rect 24 14142 260 14378
rect 12820 14142 13056 14378
rect 24 13822 260 14058
rect 12820 13822 13056 14058
rect 24 13502 260 13738
rect 12820 13502 13056 13738
rect 24 13182 260 13418
rect 12820 13182 13056 13418
rect 24 12862 260 13098
rect 12820 12862 13056 13098
rect 24 12542 260 12778
rect 12820 12542 13056 12778
rect 24 12222 260 12458
rect 12820 12222 13056 12458
rect 24 11902 260 12138
rect 12820 11902 13056 12138
rect 24 11582 260 11818
rect 12820 11582 13056 11818
rect 24 11262 260 11498
rect 12820 11262 13056 11498
rect 24 10942 260 11178
rect 12820 10942 13056 11178
rect 24 10622 260 10858
rect 12820 10622 13056 10858
rect 24 10302 260 10538
rect 12820 10302 13056 10538
rect 24 9982 260 10218
rect 12820 9982 13056 10218
rect 24 9662 260 9898
rect 12820 9662 13056 9898
rect 24 9342 260 9578
rect 12820 9342 13056 9578
rect 24 9022 260 9258
rect 12820 9022 13056 9258
rect 24 8702 260 8938
rect 12820 8702 13056 8938
rect 24 8382 260 8618
rect 12820 8382 13056 8618
rect 24 8062 260 8298
rect 12820 8200 13056 8298
rect 12820 8062 13056 8200
rect 24 7742 260 7978
rect 12820 7742 13056 7978
rect 24 7422 260 7658
rect 12820 7422 13056 7658
rect 24 7102 260 7338
rect 12820 7102 13056 7338
rect 24 6782 260 7018
rect 12820 6782 13056 7018
rect 24 6462 260 6698
rect 12820 6462 13056 6698
rect 24 6142 260 6378
rect 12820 6142 13056 6378
rect 24 5822 260 6058
rect 12820 5822 13056 6058
rect 24 5502 260 5738
rect 12820 5502 13056 5738
rect 24 5182 260 5418
rect 12820 5182 13056 5418
rect 24 4862 260 5098
rect 12820 4862 13056 5098
rect 24 4542 260 4778
rect 12820 4542 13056 4778
rect 24 4222 260 4458
rect 12820 4222 13056 4458
rect 24 3902 260 4138
rect 12820 3902 13056 4138
rect 24 3582 260 3818
rect 12820 3582 13056 3818
rect 24 3262 260 3498
rect 12820 3262 13056 3498
rect 24 2942 260 3178
rect 12820 2942 13056 3178
rect 24 2622 260 2858
rect 12820 2622 13056 2858
rect 24 2302 260 2538
rect 12820 2302 13056 2538
rect 24 1982 260 2218
rect 12820 1982 13056 2218
rect 24 1662 260 1898
rect 12820 1662 13056 1898
rect 24 1342 260 1578
rect 12820 1342 13056 1578
rect 24 1022 260 1258
rect 12820 1022 13056 1258
rect 24 702 260 938
rect 12820 702 13056 938
rect 24 382 260 618
rect 12820 382 13056 618
rect 24 24 260 260
rect 502 24 738 260
rect 822 24 1058 260
rect 1142 24 1378 260
rect 1462 24 1698 260
rect 1782 24 2018 260
rect 2102 24 2338 260
rect 2422 24 2658 260
rect 2742 24 2978 260
rect 3062 24 3298 260
rect 3382 24 3618 260
rect 3702 24 3938 260
rect 4022 24 4258 260
rect 4342 24 4578 260
rect 4662 24 4898 260
rect 4982 24 5218 260
rect 5302 24 5538 260
rect 5622 24 5858 260
rect 5942 24 6178 260
rect 6262 24 6498 260
rect 6582 24 6818 260
rect 6902 24 7138 260
rect 7222 24 7458 260
rect 7542 24 7778 260
rect 7862 24 8098 260
rect 8182 24 8418 260
rect 8502 24 8738 260
rect 8822 24 9058 260
rect 9142 24 9378 260
rect 9462 24 9698 260
rect 9782 24 10018 260
rect 10102 24 10338 260
rect 10422 24 10658 260
rect 10742 24 10978 260
rect 11062 24 11298 260
rect 11382 24 11618 260
rect 11702 24 11938 260
rect 12022 24 12258 260
rect 12342 24 12578 260
rect 12820 24 13056 260
<< metal5 >>
rect 4400 15400 8600 16200
rect 0 15056 13080 15080
rect 0 14820 24 15056
rect 260 14820 502 15056
rect 738 14820 822 15056
rect 1058 14820 1142 15056
rect 1378 14820 1462 15056
rect 1698 14820 1782 15056
rect 2018 14820 2102 15056
rect 2338 14820 2422 15056
rect 2658 14820 2742 15056
rect 2978 14820 3062 15056
rect 3298 14820 3382 15056
rect 3618 14820 3702 15056
rect 3938 14820 4022 15056
rect 4258 14820 4342 15056
rect 4578 14820 4662 15056
rect 4898 14820 4982 15056
rect 5218 14820 5302 15056
rect 5538 14820 5622 15056
rect 5858 14820 5942 15056
rect 6178 14820 6262 15056
rect 6498 14820 6582 15056
rect 6818 14820 6902 15056
rect 7138 14820 7222 15056
rect 7458 14820 7542 15056
rect 7778 14820 7862 15056
rect 8098 14820 8182 15056
rect 8418 14820 8502 15056
rect 8738 14820 8822 15056
rect 9058 14820 9142 15056
rect 9378 14820 9462 15056
rect 9698 14820 9782 15056
rect 10018 14820 10102 15056
rect 10338 14820 10422 15056
rect 10658 14820 10742 15056
rect 10978 14820 11062 15056
rect 11298 14820 11382 15056
rect 11618 14820 11702 15056
rect 11938 14820 12022 15056
rect 12258 14820 12342 15056
rect 12578 14820 12820 15056
rect 13056 14820 13080 15056
rect 0 14698 13080 14820
rect 0 14462 24 14698
rect 260 14462 12820 14698
rect 13056 14462 13080 14698
rect 0 14378 13080 14462
rect 0 14142 24 14378
rect 260 14142 12820 14378
rect 13056 14142 13080 14378
rect 0 14058 13080 14142
rect 0 13822 24 14058
rect 260 13822 12820 14058
rect 13056 13822 13080 14058
rect 0 13738 13080 13822
rect 0 13502 24 13738
rect 260 13502 12820 13738
rect 13056 13502 13080 13738
rect 0 13418 13080 13502
rect 0 13182 24 13418
rect 260 13182 12820 13418
rect 13056 13182 13080 13418
rect 0 13098 13080 13182
rect 0 12862 24 13098
rect 260 12862 12820 13098
rect 13056 12862 13080 13098
rect 0 12778 13080 12862
rect 0 12542 24 12778
rect 260 12542 12820 12778
rect 13056 12542 13080 12778
rect 0 12458 13080 12542
rect 0 12222 24 12458
rect 260 12222 12820 12458
rect 13056 12222 13080 12458
rect 0 12138 13080 12222
rect 0 11902 24 12138
rect 260 11902 12820 12138
rect 13056 11902 13080 12138
rect 0 11818 13080 11902
rect 0 11582 24 11818
rect 260 11582 12820 11818
rect 13056 11582 13080 11818
rect 0 11498 13080 11582
rect 0 11262 24 11498
rect 260 11262 12820 11498
rect 13056 11262 13080 11498
rect 0 11178 13080 11262
rect 0 10942 24 11178
rect 260 10942 12820 11178
rect 13056 10942 13080 11178
rect 0 10858 13080 10942
rect 0 10622 24 10858
rect 260 10622 12820 10858
rect 13056 10622 13080 10858
rect 0 10538 13080 10622
rect 0 10302 24 10538
rect 260 10302 12820 10538
rect 13056 10302 13080 10538
rect 0 10218 13080 10302
rect 0 9982 24 10218
rect 260 9982 12820 10218
rect 13056 9982 13080 10218
rect 0 9898 13080 9982
rect 0 9662 24 9898
rect 260 9662 12820 9898
rect 13056 9662 13080 9898
rect 0 9578 13080 9662
rect 0 9342 24 9578
rect 260 9342 12820 9578
rect 13056 9342 13080 9578
rect 0 9258 13080 9342
rect 0 9022 24 9258
rect 260 9022 12820 9258
rect 13056 9022 13080 9258
rect 0 8938 13080 9022
rect 0 8702 24 8938
rect 260 8702 12820 8938
rect 13056 8702 13080 8938
rect 0 8618 13080 8702
rect 0 8382 24 8618
rect 260 8382 12820 8618
rect 13056 8382 13080 8618
rect 0 8298 13080 8382
rect 0 8062 24 8298
rect 260 8062 12820 8298
rect 13056 8062 13080 8298
rect 0 7978 13080 8062
rect 0 7742 24 7978
rect 260 7742 12820 7978
rect 13056 7742 13080 7978
rect 0 7658 13080 7742
rect 0 7422 24 7658
rect 260 7422 12820 7658
rect 13056 7422 13080 7658
rect 0 7338 13080 7422
rect 0 7102 24 7338
rect 260 7102 12820 7338
rect 13056 7102 13080 7338
rect 0 7018 13080 7102
rect 0 6782 24 7018
rect 260 6782 12820 7018
rect 13056 6782 13080 7018
rect 0 6698 13080 6782
rect 0 6462 24 6698
rect 260 6462 12820 6698
rect 13056 6462 13080 6698
rect 0 6378 13080 6462
rect 0 6142 24 6378
rect 260 6142 12820 6378
rect 13056 6142 13080 6378
rect 0 6058 13080 6142
rect 0 5822 24 6058
rect 260 5822 12820 6058
rect 13056 5822 13080 6058
rect 0 5738 13080 5822
rect 0 5502 24 5738
rect 260 5502 12820 5738
rect 13056 5502 13080 5738
rect 0 5418 13080 5502
rect 0 5182 24 5418
rect 260 5182 12820 5418
rect 13056 5182 13080 5418
rect 0 5098 13080 5182
rect 0 4862 24 5098
rect 260 4862 12820 5098
rect 13056 4862 13080 5098
rect 0 4778 13080 4862
rect 0 4542 24 4778
rect 260 4542 12820 4778
rect 13056 4542 13080 4778
rect 0 4458 13080 4542
rect 0 4222 24 4458
rect 260 4222 12820 4458
rect 13056 4222 13080 4458
rect 0 4138 13080 4222
rect 0 3902 24 4138
rect 260 3902 12820 4138
rect 13056 3902 13080 4138
rect 0 3818 13080 3902
rect 0 3582 24 3818
rect 260 3582 12820 3818
rect 13056 3582 13080 3818
rect 0 3498 13080 3582
rect 0 3262 24 3498
rect 260 3262 12820 3498
rect 13056 3262 13080 3498
rect 0 3178 13080 3262
rect 0 2942 24 3178
rect 260 2942 12820 3178
rect 13056 2942 13080 3178
rect 0 2858 13080 2942
rect 0 2622 24 2858
rect 260 2622 12820 2858
rect 13056 2622 13080 2858
rect 0 2538 13080 2622
rect 0 2302 24 2538
rect 260 2302 12820 2538
rect 13056 2302 13080 2538
rect 0 2218 13080 2302
rect 0 1982 24 2218
rect 260 1982 12820 2218
rect 13056 1982 13080 2218
rect 0 1898 13080 1982
rect 0 1662 24 1898
rect 260 1662 12820 1898
rect 13056 1662 13080 1898
rect 0 1578 13080 1662
rect 0 1342 24 1578
rect 260 1342 12820 1578
rect 13056 1342 13080 1578
rect 0 1258 13080 1342
rect 0 1022 24 1258
rect 260 1022 12820 1258
rect 13056 1022 13080 1258
rect 0 938 13080 1022
rect 0 702 24 938
rect 260 702 12820 938
rect 13056 702 13080 938
rect 0 618 13080 702
rect 0 382 24 618
rect 260 382 12820 618
rect 13056 382 13080 618
rect 0 260 13080 382
rect 0 24 24 260
rect 260 24 502 260
rect 738 24 822 260
rect 1058 24 1142 260
rect 1378 24 1462 260
rect 1698 24 1782 260
rect 2018 24 2102 260
rect 2338 24 2422 260
rect 2658 24 2742 260
rect 2978 24 3062 260
rect 3298 24 3382 260
rect 3618 24 3702 260
rect 3938 24 4022 260
rect 4258 24 4342 260
rect 4578 24 4662 260
rect 4898 24 4982 260
rect 5218 24 5302 260
rect 5538 24 5622 260
rect 5858 24 5942 260
rect 6178 24 6262 260
rect 6498 24 6582 260
rect 6818 24 6902 260
rect 7138 24 7222 260
rect 7458 24 7542 260
rect 7778 24 7862 260
rect 8098 24 8182 260
rect 8418 24 8502 260
rect 8738 24 8822 260
rect 9058 24 9142 260
rect 9378 24 9462 260
rect 9698 24 9782 260
rect 10018 24 10102 260
rect 10338 24 10422 260
rect 10658 24 10742 260
rect 10978 24 11062 260
rect 11298 24 11382 260
rect 11618 24 11702 260
rect 11938 24 12022 260
rect 12258 24 12342 260
rect 12578 24 12820 260
rect 13056 24 13080 260
rect 0 0 13080 24
<< glass >>
rect 540 540 12540 14540
<< labels >>
flabel metal5 4400 15400 8600 16200 0 FreeSans 6400 0 0 0 pad
port 1 nsew
flabel metal1 1700 1600 2160 2200 0 FreeSans 3200 0 0 0 GND
flabel metal5 s 260 260 12820 14820 0 FreeSans 2000 0 0 0 PAD
<< end >>
