magic
tech sky130A
magscale 1 2
timestamp 1717597427
<< error_p >>
rect 1982 29160 2302 29230
rect 366 28916 606 28940
rect 366 28724 390 28916
rect 582 28724 606 28916
rect 1982 28920 2006 29160
rect 2232 28920 2246 29160
rect 2256 28920 2302 29160
rect 5982 29160 6302 29230
rect 1982 28896 2302 28920
rect 4366 28916 4606 28940
rect 366 28700 606 28724
rect 4366 28724 4390 28916
rect 4582 28724 4606 28916
rect 5982 28920 6006 29160
rect 6232 28920 6246 29160
rect 6256 28920 6302 29160
rect 9982 29160 10302 29230
rect 5982 28896 6302 28920
rect 8366 28916 8606 28940
rect 2852 28709 2996 28714
rect 2852 28639 2857 28709
rect 2991 28639 2996 28709
rect 4366 28700 4606 28724
rect 8366 28724 8390 28916
rect 8582 28724 8606 28916
rect 9982 28920 10006 29160
rect 10232 28920 10246 29160
rect 10256 28920 10302 29160
rect 13982 29160 14302 29230
rect 9982 28896 10302 28920
rect 12366 28916 12606 28940
rect 6852 28709 6996 28714
rect 2852 28634 2996 28639
rect 6852 28639 6857 28709
rect 6991 28639 6996 28709
rect 8366 28700 8606 28724
rect 12366 28724 12390 28916
rect 12582 28724 12606 28916
rect 13982 28920 14006 29160
rect 14232 28920 14246 29160
rect 14256 28920 14302 29160
rect 17982 29160 18302 29230
rect 13982 28896 14302 28920
rect 16366 28916 16606 28940
rect 10852 28709 10996 28714
rect 6852 28634 6996 28639
rect 10852 28639 10857 28709
rect 10991 28639 10996 28709
rect 12366 28700 12606 28724
rect 16366 28724 16390 28916
rect 16582 28724 16606 28916
rect 17982 28920 18006 29160
rect 18232 28920 18246 29160
rect 18256 28920 18302 29160
rect 21982 29160 22302 29230
rect 17982 28896 18302 28920
rect 20366 28916 20606 28940
rect 14852 28709 14996 28714
rect 10852 28634 10996 28639
rect 14852 28639 14857 28709
rect 14991 28639 14996 28709
rect 16366 28700 16606 28724
rect 20366 28724 20390 28916
rect 20582 28724 20606 28916
rect 21982 28920 22006 29160
rect 22232 28920 22246 29160
rect 22256 28920 22302 29160
rect 25982 29160 26302 29230
rect 21982 28896 22302 28920
rect 24366 28916 24606 28940
rect 18852 28709 18996 28714
rect 14852 28634 14996 28639
rect 18852 28639 18857 28709
rect 18991 28639 18996 28709
rect 20366 28700 20606 28724
rect 24366 28724 24390 28916
rect 24582 28724 24606 28916
rect 25982 28920 26006 29160
rect 26232 28920 26246 29160
rect 26256 28920 26302 29160
rect 29982 29160 30302 29230
rect 25982 28896 26302 28920
rect 28366 28916 28606 28940
rect 22852 28709 22996 28714
rect 18852 28634 18996 28639
rect 22852 28639 22857 28709
rect 22991 28639 22996 28709
rect 24366 28700 24606 28724
rect 28366 28724 28390 28916
rect 28582 28724 28606 28916
rect 29982 28920 30006 29160
rect 30232 28920 30246 29160
rect 30256 28920 30302 29160
rect 33982 29160 34302 29230
rect 29982 28896 30302 28920
rect 32366 28916 32606 28940
rect 26852 28709 26996 28714
rect 22852 28634 22996 28639
rect 26852 28639 26857 28709
rect 26991 28639 26996 28709
rect 28366 28700 28606 28724
rect 32366 28724 32390 28916
rect 32582 28724 32606 28916
rect 33982 28920 34006 29160
rect 34232 28920 34246 29160
rect 34256 28920 34302 29160
rect 37982 29160 38302 29230
rect 33982 28896 34302 28920
rect 36366 28916 36606 28940
rect 30852 28709 30996 28714
rect 26852 28634 26996 28639
rect 30852 28639 30857 28709
rect 30991 28639 30996 28709
rect 32366 28700 32606 28724
rect 36366 28724 36390 28916
rect 36582 28724 36606 28916
rect 37982 28920 38006 29160
rect 38232 28920 38246 29160
rect 38256 28920 38302 29160
rect 37982 28896 38302 28920
rect 34852 28709 34996 28714
rect 30852 28634 30996 28639
rect 34852 28639 34857 28709
rect 34991 28639 34996 28709
rect 36366 28700 36606 28724
rect 38852 28709 38996 28714
rect 34852 28634 34996 28639
rect 38852 28639 38857 28709
rect 38991 28639 38996 28709
rect 38852 28634 38996 28639
rect 2366 28559 2546 28560
rect 2366 28381 2367 28559
rect 2545 28381 2546 28559
rect 2366 28380 2546 28381
rect 6366 28559 6546 28560
rect 6366 28381 6367 28559
rect 6545 28381 6546 28559
rect 6366 28380 6546 28381
rect 10366 28559 10546 28560
rect 10366 28381 10367 28559
rect 10545 28381 10546 28559
rect 10366 28380 10546 28381
rect 14366 28559 14546 28560
rect 14366 28381 14367 28559
rect 14545 28381 14546 28559
rect 14366 28380 14546 28381
rect 18366 28559 18546 28560
rect 18366 28381 18367 28559
rect 18545 28381 18546 28559
rect 18366 28380 18546 28381
rect 22366 28559 22546 28560
rect 22366 28381 22367 28559
rect 22545 28381 22546 28559
rect 22366 28380 22546 28381
rect 26366 28559 26546 28560
rect 26366 28381 26367 28559
rect 26545 28381 26546 28559
rect 26366 28380 26546 28381
rect 30366 28559 30546 28560
rect 30366 28381 30367 28559
rect 30545 28381 30546 28559
rect 30366 28380 30546 28381
rect 34366 28559 34546 28560
rect 34366 28381 34367 28559
rect 34545 28381 34546 28559
rect 34366 28380 34546 28381
rect 38366 28559 38546 28560
rect 38366 28381 38367 28559
rect 38545 28381 38546 28559
rect 38366 28380 38546 28381
rect 366 28039 546 28040
rect 366 27861 367 28039
rect 545 27861 546 28039
rect 4366 28039 4546 28040
rect 3734 27984 3740 27990
rect 3780 27984 3786 27990
rect 3728 27978 3734 27984
rect 3786 27978 3792 27984
rect 3728 27928 3734 27934
rect 3786 27928 3792 27934
rect 3734 27922 3740 27928
rect 3780 27922 3786 27928
rect 366 27860 546 27861
rect 4366 27861 4367 28039
rect 4545 27861 4546 28039
rect 8366 28039 8546 28040
rect 7734 27984 7740 27990
rect 7780 27984 7786 27990
rect 7728 27978 7734 27984
rect 7786 27978 7792 27984
rect 7728 27928 7734 27934
rect 7786 27928 7792 27934
rect 7734 27922 7740 27928
rect 7780 27922 7786 27928
rect 4366 27860 4546 27861
rect 8366 27861 8367 28039
rect 8545 27861 8546 28039
rect 12366 28039 12546 28040
rect 11734 27984 11740 27990
rect 11780 27984 11786 27990
rect 11728 27978 11734 27984
rect 11786 27978 11792 27984
rect 11728 27928 11734 27934
rect 11786 27928 11792 27934
rect 11734 27922 11740 27928
rect 11780 27922 11786 27928
rect 8366 27860 8546 27861
rect 12366 27861 12367 28039
rect 12545 27861 12546 28039
rect 16366 28039 16546 28040
rect 15734 27984 15740 27990
rect 15780 27984 15786 27990
rect 15728 27978 15734 27984
rect 15786 27978 15792 27984
rect 15728 27928 15734 27934
rect 15786 27928 15792 27934
rect 15734 27922 15740 27928
rect 15780 27922 15786 27928
rect 12366 27860 12546 27861
rect 16366 27861 16367 28039
rect 16545 27861 16546 28039
rect 20366 28039 20546 28040
rect 19734 27984 19740 27990
rect 19780 27984 19786 27990
rect 19728 27978 19734 27984
rect 19786 27978 19792 27984
rect 19728 27928 19734 27934
rect 19786 27928 19792 27934
rect 19734 27922 19740 27928
rect 19780 27922 19786 27928
rect 16366 27860 16546 27861
rect 20366 27861 20367 28039
rect 20545 27861 20546 28039
rect 24366 28039 24546 28040
rect 23734 27984 23740 27990
rect 23780 27984 23786 27990
rect 23728 27978 23734 27984
rect 23786 27978 23792 27984
rect 23728 27928 23734 27934
rect 23786 27928 23792 27934
rect 23734 27922 23740 27928
rect 23780 27922 23786 27928
rect 20366 27860 20546 27861
rect 24366 27861 24367 28039
rect 24545 27861 24546 28039
rect 28366 28039 28546 28040
rect 27734 27984 27740 27990
rect 27780 27984 27786 27990
rect 27728 27978 27734 27984
rect 27786 27978 27792 27984
rect 27728 27928 27734 27934
rect 27786 27928 27792 27934
rect 27734 27922 27740 27928
rect 27780 27922 27786 27928
rect 24366 27860 24546 27861
rect 28366 27861 28367 28039
rect 28545 27861 28546 28039
rect 32366 28039 32546 28040
rect 31734 27984 31740 27990
rect 31780 27984 31786 27990
rect 31728 27978 31734 27984
rect 31786 27978 31792 27984
rect 31728 27928 31734 27934
rect 31786 27928 31792 27934
rect 31734 27922 31740 27928
rect 31780 27922 31786 27928
rect 28366 27860 28546 27861
rect 32366 27861 32367 28039
rect 32545 27861 32546 28039
rect 36366 28039 36546 28040
rect 35734 27984 35740 27990
rect 35780 27984 35786 27990
rect 35728 27978 35734 27984
rect 35786 27978 35792 27984
rect 35728 27928 35734 27934
rect 35786 27928 35792 27934
rect 35734 27922 35740 27928
rect 35780 27922 35786 27928
rect 32366 27860 32546 27861
rect 36366 27861 36367 28039
rect 36545 27861 36546 28039
rect 39734 27984 39740 27990
rect 39780 27984 39786 27990
rect 39728 27978 39734 27984
rect 39786 27978 39792 27984
rect 39728 27928 39734 27934
rect 39786 27928 39792 27934
rect 39734 27922 39740 27928
rect 39780 27922 39786 27928
rect 36366 27860 36546 27861
rect 3262 27808 3268 27814
rect 3308 27808 3314 27814
rect 7262 27808 7268 27814
rect 7308 27808 7314 27814
rect 11262 27808 11268 27814
rect 11308 27808 11314 27814
rect 15262 27808 15268 27814
rect 15308 27808 15314 27814
rect 19262 27808 19268 27814
rect 19308 27808 19314 27814
rect 23262 27808 23268 27814
rect 23308 27808 23314 27814
rect 27262 27808 27268 27814
rect 27308 27808 27314 27814
rect 31262 27808 31268 27814
rect 31308 27808 31314 27814
rect 35262 27808 35268 27814
rect 35308 27808 35314 27814
rect 39262 27808 39268 27814
rect 39308 27808 39314 27814
rect 3256 27802 3262 27808
rect 3314 27802 3320 27808
rect 7256 27802 7262 27808
rect 7314 27802 7320 27808
rect 11256 27802 11262 27808
rect 11314 27802 11320 27808
rect 15256 27802 15262 27808
rect 15314 27802 15320 27808
rect 19256 27802 19262 27808
rect 19314 27802 19320 27808
rect 23256 27802 23262 27808
rect 23314 27802 23320 27808
rect 27256 27802 27262 27808
rect 27314 27802 27320 27808
rect 31256 27802 31262 27808
rect 31314 27802 31320 27808
rect 35256 27802 35262 27808
rect 35314 27802 35320 27808
rect 39256 27802 39262 27808
rect 39314 27802 39320 27808
rect 3256 27756 3262 27762
rect 3314 27756 3320 27762
rect 7256 27756 7262 27762
rect 7314 27756 7320 27762
rect 11256 27756 11262 27762
rect 11314 27756 11320 27762
rect 15256 27756 15262 27762
rect 15314 27756 15320 27762
rect 19256 27756 19262 27762
rect 19314 27756 19320 27762
rect 23256 27756 23262 27762
rect 23314 27756 23320 27762
rect 27256 27756 27262 27762
rect 27314 27756 27320 27762
rect 31256 27756 31262 27762
rect 31314 27756 31320 27762
rect 35256 27756 35262 27762
rect 35314 27756 35320 27762
rect 39256 27756 39262 27762
rect 39314 27756 39320 27762
rect 3262 27750 3268 27756
rect 3308 27750 3314 27756
rect 7262 27750 7268 27756
rect 7308 27750 7314 27756
rect 11262 27750 11268 27756
rect 11308 27750 11314 27756
rect 15262 27750 15268 27756
rect 15308 27750 15314 27756
rect 19262 27750 19268 27756
rect 19308 27750 19314 27756
rect 23262 27750 23268 27756
rect 23308 27750 23314 27756
rect 27262 27750 27268 27756
rect 27308 27750 27314 27756
rect 31262 27750 31268 27756
rect 31308 27750 31314 27756
rect 35262 27750 35268 27756
rect 35308 27750 35314 27756
rect 39262 27750 39268 27756
rect 39308 27750 39314 27756
rect 2386 27296 2626 27320
rect 2386 27104 2410 27296
rect 2602 27104 2626 27296
rect 2386 27080 2626 27104
rect 6386 27296 6626 27320
rect 6386 27104 6410 27296
rect 6602 27104 6626 27296
rect 6386 27080 6626 27104
rect 10386 27296 10626 27320
rect 10386 27104 10410 27296
rect 10602 27104 10626 27296
rect 10386 27080 10626 27104
rect 14386 27296 14626 27320
rect 14386 27104 14410 27296
rect 14602 27104 14626 27296
rect 14386 27080 14626 27104
rect 18386 27296 18626 27320
rect 18386 27104 18410 27296
rect 18602 27104 18626 27296
rect 18386 27080 18626 27104
rect 22386 27296 22626 27320
rect 22386 27104 22410 27296
rect 22602 27104 22626 27296
rect 22386 27080 22626 27104
rect 26386 27296 26626 27320
rect 26386 27104 26410 27296
rect 26602 27104 26626 27296
rect 26386 27080 26626 27104
rect 30386 27296 30626 27320
rect 30386 27104 30410 27296
rect 30602 27104 30626 27296
rect 30386 27080 30626 27104
rect 34386 27296 34626 27320
rect 34386 27104 34410 27296
rect 34602 27104 34626 27296
rect 34386 27080 34626 27104
rect 38386 27296 38626 27320
rect 38386 27104 38410 27296
rect 38602 27104 38626 27296
rect 38386 27080 38626 27104
rect 1982 26160 2302 26230
rect 366 25916 606 25940
rect 366 25724 390 25916
rect 582 25724 606 25916
rect 1982 25920 2006 26160
rect 2232 25920 2246 26160
rect 2256 25920 2302 26160
rect 5982 26160 6302 26230
rect 1982 25896 2302 25920
rect 4366 25916 4606 25940
rect 366 25700 606 25724
rect 4366 25724 4390 25916
rect 4582 25724 4606 25916
rect 5982 25920 6006 26160
rect 6232 25920 6246 26160
rect 6256 25920 6302 26160
rect 9982 26160 10302 26230
rect 5982 25896 6302 25920
rect 8366 25916 8606 25940
rect 2852 25709 2996 25714
rect 2852 25639 2857 25709
rect 2991 25639 2996 25709
rect 4366 25700 4606 25724
rect 8366 25724 8390 25916
rect 8582 25724 8606 25916
rect 9982 25920 10006 26160
rect 10232 25920 10246 26160
rect 10256 25920 10302 26160
rect 13982 26160 14302 26230
rect 9982 25896 10302 25920
rect 12366 25916 12606 25940
rect 6852 25709 6996 25714
rect 2852 25634 2996 25639
rect 6852 25639 6857 25709
rect 6991 25639 6996 25709
rect 8366 25700 8606 25724
rect 12366 25724 12390 25916
rect 12582 25724 12606 25916
rect 13982 25920 14006 26160
rect 14232 25920 14246 26160
rect 14256 25920 14302 26160
rect 17982 26160 18302 26230
rect 13982 25896 14302 25920
rect 16366 25916 16606 25940
rect 10852 25709 10996 25714
rect 6852 25634 6996 25639
rect 10852 25639 10857 25709
rect 10991 25639 10996 25709
rect 12366 25700 12606 25724
rect 16366 25724 16390 25916
rect 16582 25724 16606 25916
rect 17982 25920 18006 26160
rect 18232 25920 18246 26160
rect 18256 25920 18302 26160
rect 21982 26160 22302 26230
rect 17982 25896 18302 25920
rect 20366 25916 20606 25940
rect 14852 25709 14996 25714
rect 10852 25634 10996 25639
rect 14852 25639 14857 25709
rect 14991 25639 14996 25709
rect 16366 25700 16606 25724
rect 20366 25724 20390 25916
rect 20582 25724 20606 25916
rect 21982 25920 22006 26160
rect 22232 25920 22246 26160
rect 22256 25920 22302 26160
rect 25982 26160 26302 26230
rect 21982 25896 22302 25920
rect 24366 25916 24606 25940
rect 18852 25709 18996 25714
rect 14852 25634 14996 25639
rect 18852 25639 18857 25709
rect 18991 25639 18996 25709
rect 20366 25700 20606 25724
rect 24366 25724 24390 25916
rect 24582 25724 24606 25916
rect 25982 25920 26006 26160
rect 26232 25920 26246 26160
rect 26256 25920 26302 26160
rect 29982 26160 30302 26230
rect 25982 25896 26302 25920
rect 28366 25916 28606 25940
rect 22852 25709 22996 25714
rect 18852 25634 18996 25639
rect 22852 25639 22857 25709
rect 22991 25639 22996 25709
rect 24366 25700 24606 25724
rect 28366 25724 28390 25916
rect 28582 25724 28606 25916
rect 29982 25920 30006 26160
rect 30232 25920 30246 26160
rect 30256 25920 30302 26160
rect 33982 26160 34302 26230
rect 29982 25896 30302 25920
rect 32366 25916 32606 25940
rect 26852 25709 26996 25714
rect 22852 25634 22996 25639
rect 26852 25639 26857 25709
rect 26991 25639 26996 25709
rect 28366 25700 28606 25724
rect 32366 25724 32390 25916
rect 32582 25724 32606 25916
rect 33982 25920 34006 26160
rect 34232 25920 34246 26160
rect 34256 25920 34302 26160
rect 37982 26160 38302 26230
rect 33982 25896 34302 25920
rect 36366 25916 36606 25940
rect 30852 25709 30996 25714
rect 26852 25634 26996 25639
rect 30852 25639 30857 25709
rect 30991 25639 30996 25709
rect 32366 25700 32606 25724
rect 36366 25724 36390 25916
rect 36582 25724 36606 25916
rect 37982 25920 38006 26160
rect 38232 25920 38246 26160
rect 38256 25920 38302 26160
rect 37982 25896 38302 25920
rect 34852 25709 34996 25714
rect 30852 25634 30996 25639
rect 34852 25639 34857 25709
rect 34991 25639 34996 25709
rect 36366 25700 36606 25724
rect 38852 25709 38996 25714
rect 34852 25634 34996 25639
rect 38852 25639 38857 25709
rect 38991 25639 38996 25709
rect 38852 25634 38996 25639
rect 2366 25559 2546 25560
rect 2366 25381 2367 25559
rect 2545 25381 2546 25559
rect 2366 25380 2546 25381
rect 6366 25559 6546 25560
rect 6366 25381 6367 25559
rect 6545 25381 6546 25559
rect 6366 25380 6546 25381
rect 10366 25559 10546 25560
rect 10366 25381 10367 25559
rect 10545 25381 10546 25559
rect 10366 25380 10546 25381
rect 14366 25559 14546 25560
rect 14366 25381 14367 25559
rect 14545 25381 14546 25559
rect 14366 25380 14546 25381
rect 18366 25559 18546 25560
rect 18366 25381 18367 25559
rect 18545 25381 18546 25559
rect 18366 25380 18546 25381
rect 22366 25559 22546 25560
rect 22366 25381 22367 25559
rect 22545 25381 22546 25559
rect 22366 25380 22546 25381
rect 26366 25559 26546 25560
rect 26366 25381 26367 25559
rect 26545 25381 26546 25559
rect 26366 25380 26546 25381
rect 30366 25559 30546 25560
rect 30366 25381 30367 25559
rect 30545 25381 30546 25559
rect 30366 25380 30546 25381
rect 34366 25559 34546 25560
rect 34366 25381 34367 25559
rect 34545 25381 34546 25559
rect 34366 25380 34546 25381
rect 38366 25559 38546 25560
rect 38366 25381 38367 25559
rect 38545 25381 38546 25559
rect 38366 25380 38546 25381
rect 366 25039 546 25040
rect 366 24861 367 25039
rect 545 24861 546 25039
rect 4366 25039 4546 25040
rect 3734 24984 3740 24990
rect 3780 24984 3786 24990
rect 3728 24978 3734 24984
rect 3786 24978 3792 24984
rect 3728 24928 3734 24934
rect 3786 24928 3792 24934
rect 3734 24922 3740 24928
rect 3780 24922 3786 24928
rect 366 24860 546 24861
rect 4366 24861 4367 25039
rect 4545 24861 4546 25039
rect 8366 25039 8546 25040
rect 7734 24984 7740 24990
rect 7780 24984 7786 24990
rect 7728 24978 7734 24984
rect 7786 24978 7792 24984
rect 7728 24928 7734 24934
rect 7786 24928 7792 24934
rect 7734 24922 7740 24928
rect 7780 24922 7786 24928
rect 4366 24860 4546 24861
rect 8366 24861 8367 25039
rect 8545 24861 8546 25039
rect 12366 25039 12546 25040
rect 11734 24984 11740 24990
rect 11780 24984 11786 24990
rect 11728 24978 11734 24984
rect 11786 24978 11792 24984
rect 11728 24928 11734 24934
rect 11786 24928 11792 24934
rect 11734 24922 11740 24928
rect 11780 24922 11786 24928
rect 8366 24860 8546 24861
rect 12366 24861 12367 25039
rect 12545 24861 12546 25039
rect 16366 25039 16546 25040
rect 15734 24984 15740 24990
rect 15780 24984 15786 24990
rect 15728 24978 15734 24984
rect 15786 24978 15792 24984
rect 15728 24928 15734 24934
rect 15786 24928 15792 24934
rect 15734 24922 15740 24928
rect 15780 24922 15786 24928
rect 12366 24860 12546 24861
rect 16366 24861 16367 25039
rect 16545 24861 16546 25039
rect 20366 25039 20546 25040
rect 19734 24984 19740 24990
rect 19780 24984 19786 24990
rect 19728 24978 19734 24984
rect 19786 24978 19792 24984
rect 19728 24928 19734 24934
rect 19786 24928 19792 24934
rect 19734 24922 19740 24928
rect 19780 24922 19786 24928
rect 16366 24860 16546 24861
rect 20366 24861 20367 25039
rect 20545 24861 20546 25039
rect 24366 25039 24546 25040
rect 23734 24984 23740 24990
rect 23780 24984 23786 24990
rect 23728 24978 23734 24984
rect 23786 24978 23792 24984
rect 23728 24928 23734 24934
rect 23786 24928 23792 24934
rect 23734 24922 23740 24928
rect 23780 24922 23786 24928
rect 20366 24860 20546 24861
rect 24366 24861 24367 25039
rect 24545 24861 24546 25039
rect 28366 25039 28546 25040
rect 27734 24984 27740 24990
rect 27780 24984 27786 24990
rect 27728 24978 27734 24984
rect 27786 24978 27792 24984
rect 27728 24928 27734 24934
rect 27786 24928 27792 24934
rect 27734 24922 27740 24928
rect 27780 24922 27786 24928
rect 24366 24860 24546 24861
rect 28366 24861 28367 25039
rect 28545 24861 28546 25039
rect 32366 25039 32546 25040
rect 31734 24984 31740 24990
rect 31780 24984 31786 24990
rect 31728 24978 31734 24984
rect 31786 24978 31792 24984
rect 31728 24928 31734 24934
rect 31786 24928 31792 24934
rect 31734 24922 31740 24928
rect 31780 24922 31786 24928
rect 28366 24860 28546 24861
rect 32366 24861 32367 25039
rect 32545 24861 32546 25039
rect 36366 25039 36546 25040
rect 35734 24984 35740 24990
rect 35780 24984 35786 24990
rect 35728 24978 35734 24984
rect 35786 24978 35792 24984
rect 35728 24928 35734 24934
rect 35786 24928 35792 24934
rect 35734 24922 35740 24928
rect 35780 24922 35786 24928
rect 32366 24860 32546 24861
rect 36366 24861 36367 25039
rect 36545 24861 36546 25039
rect 39734 24984 39740 24990
rect 39780 24984 39786 24990
rect 39728 24978 39734 24984
rect 39786 24978 39792 24984
rect 39728 24928 39734 24934
rect 39786 24928 39792 24934
rect 39734 24922 39740 24928
rect 39780 24922 39786 24928
rect 36366 24860 36546 24861
rect 3262 24808 3268 24814
rect 3308 24808 3314 24814
rect 7262 24808 7268 24814
rect 7308 24808 7314 24814
rect 11262 24808 11268 24814
rect 11308 24808 11314 24814
rect 15262 24808 15268 24814
rect 15308 24808 15314 24814
rect 19262 24808 19268 24814
rect 19308 24808 19314 24814
rect 23262 24808 23268 24814
rect 23308 24808 23314 24814
rect 27262 24808 27268 24814
rect 27308 24808 27314 24814
rect 31262 24808 31268 24814
rect 31308 24808 31314 24814
rect 35262 24808 35268 24814
rect 35308 24808 35314 24814
rect 39262 24808 39268 24814
rect 39308 24808 39314 24814
rect 3256 24802 3262 24808
rect 3314 24802 3320 24808
rect 7256 24802 7262 24808
rect 7314 24802 7320 24808
rect 11256 24802 11262 24808
rect 11314 24802 11320 24808
rect 15256 24802 15262 24808
rect 15314 24802 15320 24808
rect 19256 24802 19262 24808
rect 19314 24802 19320 24808
rect 23256 24802 23262 24808
rect 23314 24802 23320 24808
rect 27256 24802 27262 24808
rect 27314 24802 27320 24808
rect 31256 24802 31262 24808
rect 31314 24802 31320 24808
rect 35256 24802 35262 24808
rect 35314 24802 35320 24808
rect 39256 24802 39262 24808
rect 39314 24802 39320 24808
rect 3256 24756 3262 24762
rect 3314 24756 3320 24762
rect 7256 24756 7262 24762
rect 7314 24756 7320 24762
rect 11256 24756 11262 24762
rect 11314 24756 11320 24762
rect 15256 24756 15262 24762
rect 15314 24756 15320 24762
rect 19256 24756 19262 24762
rect 19314 24756 19320 24762
rect 23256 24756 23262 24762
rect 23314 24756 23320 24762
rect 27256 24756 27262 24762
rect 27314 24756 27320 24762
rect 31256 24756 31262 24762
rect 31314 24756 31320 24762
rect 35256 24756 35262 24762
rect 35314 24756 35320 24762
rect 39256 24756 39262 24762
rect 39314 24756 39320 24762
rect 3262 24750 3268 24756
rect 3308 24750 3314 24756
rect 7262 24750 7268 24756
rect 7308 24750 7314 24756
rect 11262 24750 11268 24756
rect 11308 24750 11314 24756
rect 15262 24750 15268 24756
rect 15308 24750 15314 24756
rect 19262 24750 19268 24756
rect 19308 24750 19314 24756
rect 23262 24750 23268 24756
rect 23308 24750 23314 24756
rect 27262 24750 27268 24756
rect 27308 24750 27314 24756
rect 31262 24750 31268 24756
rect 31308 24750 31314 24756
rect 35262 24750 35268 24756
rect 35308 24750 35314 24756
rect 39262 24750 39268 24756
rect 39308 24750 39314 24756
rect 2386 24296 2626 24320
rect 2386 24104 2410 24296
rect 2602 24104 2626 24296
rect 2386 24080 2626 24104
rect 6386 24296 6626 24320
rect 6386 24104 6410 24296
rect 6602 24104 6626 24296
rect 6386 24080 6626 24104
rect 10386 24296 10626 24320
rect 10386 24104 10410 24296
rect 10602 24104 10626 24296
rect 10386 24080 10626 24104
rect 14386 24296 14626 24320
rect 14386 24104 14410 24296
rect 14602 24104 14626 24296
rect 14386 24080 14626 24104
rect 18386 24296 18626 24320
rect 18386 24104 18410 24296
rect 18602 24104 18626 24296
rect 18386 24080 18626 24104
rect 22386 24296 22626 24320
rect 22386 24104 22410 24296
rect 22602 24104 22626 24296
rect 22386 24080 22626 24104
rect 26386 24296 26626 24320
rect 26386 24104 26410 24296
rect 26602 24104 26626 24296
rect 26386 24080 26626 24104
rect 30386 24296 30626 24320
rect 30386 24104 30410 24296
rect 30602 24104 30626 24296
rect 30386 24080 30626 24104
rect 34386 24296 34626 24320
rect 34386 24104 34410 24296
rect 34602 24104 34626 24296
rect 34386 24080 34626 24104
rect 38386 24296 38626 24320
rect 38386 24104 38410 24296
rect 38602 24104 38626 24296
rect 38386 24080 38626 24104
rect 1982 23160 2302 23230
rect 366 22916 606 22940
rect 366 22724 390 22916
rect 582 22724 606 22916
rect 1982 22920 2006 23160
rect 2232 22920 2246 23160
rect 2256 22920 2302 23160
rect 5982 23160 6302 23230
rect 1982 22896 2302 22920
rect 4366 22916 4606 22940
rect 366 22700 606 22724
rect 4366 22724 4390 22916
rect 4582 22724 4606 22916
rect 5982 22920 6006 23160
rect 6232 22920 6246 23160
rect 6256 22920 6302 23160
rect 9982 23160 10302 23230
rect 5982 22896 6302 22920
rect 8366 22916 8606 22940
rect 2852 22709 2996 22714
rect 2852 22639 2857 22709
rect 2991 22639 2996 22709
rect 4366 22700 4606 22724
rect 8366 22724 8390 22916
rect 8582 22724 8606 22916
rect 9982 22920 10006 23160
rect 10232 22920 10246 23160
rect 10256 22920 10302 23160
rect 13982 23160 14302 23230
rect 9982 22896 10302 22920
rect 12366 22916 12606 22940
rect 6852 22709 6996 22714
rect 2852 22634 2996 22639
rect 6852 22639 6857 22709
rect 6991 22639 6996 22709
rect 8366 22700 8606 22724
rect 12366 22724 12390 22916
rect 12582 22724 12606 22916
rect 13982 22920 14006 23160
rect 14232 22920 14246 23160
rect 14256 22920 14302 23160
rect 17982 23160 18302 23230
rect 13982 22896 14302 22920
rect 16366 22916 16606 22940
rect 10852 22709 10996 22714
rect 6852 22634 6996 22639
rect 10852 22639 10857 22709
rect 10991 22639 10996 22709
rect 12366 22700 12606 22724
rect 16366 22724 16390 22916
rect 16582 22724 16606 22916
rect 17982 22920 18006 23160
rect 18232 22920 18246 23160
rect 18256 22920 18302 23160
rect 21982 23160 22302 23230
rect 17982 22896 18302 22920
rect 20366 22916 20606 22940
rect 14852 22709 14996 22714
rect 10852 22634 10996 22639
rect 14852 22639 14857 22709
rect 14991 22639 14996 22709
rect 16366 22700 16606 22724
rect 20366 22724 20390 22916
rect 20582 22724 20606 22916
rect 21982 22920 22006 23160
rect 22232 22920 22246 23160
rect 22256 22920 22302 23160
rect 25982 23160 26302 23230
rect 21982 22896 22302 22920
rect 24366 22916 24606 22940
rect 18852 22709 18996 22714
rect 14852 22634 14996 22639
rect 18852 22639 18857 22709
rect 18991 22639 18996 22709
rect 20366 22700 20606 22724
rect 24366 22724 24390 22916
rect 24582 22724 24606 22916
rect 25982 22920 26006 23160
rect 26232 22920 26246 23160
rect 26256 22920 26302 23160
rect 29982 23160 30302 23230
rect 25982 22896 26302 22920
rect 28366 22916 28606 22940
rect 22852 22709 22996 22714
rect 18852 22634 18996 22639
rect 22852 22639 22857 22709
rect 22991 22639 22996 22709
rect 24366 22700 24606 22724
rect 28366 22724 28390 22916
rect 28582 22724 28606 22916
rect 29982 22920 30006 23160
rect 30232 22920 30246 23160
rect 30256 22920 30302 23160
rect 33982 23160 34302 23230
rect 29982 22896 30302 22920
rect 32366 22916 32606 22940
rect 26852 22709 26996 22714
rect 22852 22634 22996 22639
rect 26852 22639 26857 22709
rect 26991 22639 26996 22709
rect 28366 22700 28606 22724
rect 32366 22724 32390 22916
rect 32582 22724 32606 22916
rect 33982 22920 34006 23160
rect 34232 22920 34246 23160
rect 34256 22920 34302 23160
rect 37982 23160 38302 23230
rect 33982 22896 34302 22920
rect 36366 22916 36606 22940
rect 30852 22709 30996 22714
rect 26852 22634 26996 22639
rect 30852 22639 30857 22709
rect 30991 22639 30996 22709
rect 32366 22700 32606 22724
rect 36366 22724 36390 22916
rect 36582 22724 36606 22916
rect 37982 22920 38006 23160
rect 38232 22920 38246 23160
rect 38256 22920 38302 23160
rect 37982 22896 38302 22920
rect 34852 22709 34996 22714
rect 30852 22634 30996 22639
rect 34852 22639 34857 22709
rect 34991 22639 34996 22709
rect 36366 22700 36606 22724
rect 38852 22709 38996 22714
rect 34852 22634 34996 22639
rect 38852 22639 38857 22709
rect 38991 22639 38996 22709
rect 38852 22634 38996 22639
rect 2366 22559 2546 22560
rect 2366 22381 2367 22559
rect 2545 22381 2546 22559
rect 2366 22380 2546 22381
rect 6366 22559 6546 22560
rect 6366 22381 6367 22559
rect 6545 22381 6546 22559
rect 6366 22380 6546 22381
rect 10366 22559 10546 22560
rect 10366 22381 10367 22559
rect 10545 22381 10546 22559
rect 10366 22380 10546 22381
rect 14366 22559 14546 22560
rect 14366 22381 14367 22559
rect 14545 22381 14546 22559
rect 14366 22380 14546 22381
rect 18366 22559 18546 22560
rect 18366 22381 18367 22559
rect 18545 22381 18546 22559
rect 18366 22380 18546 22381
rect 22366 22559 22546 22560
rect 22366 22381 22367 22559
rect 22545 22381 22546 22559
rect 22366 22380 22546 22381
rect 26366 22559 26546 22560
rect 26366 22381 26367 22559
rect 26545 22381 26546 22559
rect 26366 22380 26546 22381
rect 30366 22559 30546 22560
rect 30366 22381 30367 22559
rect 30545 22381 30546 22559
rect 30366 22380 30546 22381
rect 34366 22559 34546 22560
rect 34366 22381 34367 22559
rect 34545 22381 34546 22559
rect 34366 22380 34546 22381
rect 38366 22559 38546 22560
rect 38366 22381 38367 22559
rect 38545 22381 38546 22559
rect 38366 22380 38546 22381
rect 366 22039 546 22040
rect 366 21861 367 22039
rect 545 21861 546 22039
rect 4366 22039 4546 22040
rect 3734 21984 3740 21990
rect 3780 21984 3786 21990
rect 3728 21978 3734 21984
rect 3786 21978 3792 21984
rect 3728 21928 3734 21934
rect 3786 21928 3792 21934
rect 3734 21922 3740 21928
rect 3780 21922 3786 21928
rect 366 21860 546 21861
rect 4366 21861 4367 22039
rect 4545 21861 4546 22039
rect 8366 22039 8546 22040
rect 7734 21984 7740 21990
rect 7780 21984 7786 21990
rect 7728 21978 7734 21984
rect 7786 21978 7792 21984
rect 7728 21928 7734 21934
rect 7786 21928 7792 21934
rect 7734 21922 7740 21928
rect 7780 21922 7786 21928
rect 4366 21860 4546 21861
rect 8366 21861 8367 22039
rect 8545 21861 8546 22039
rect 12366 22039 12546 22040
rect 11734 21984 11740 21990
rect 11780 21984 11786 21990
rect 11728 21978 11734 21984
rect 11786 21978 11792 21984
rect 11728 21928 11734 21934
rect 11786 21928 11792 21934
rect 11734 21922 11740 21928
rect 11780 21922 11786 21928
rect 8366 21860 8546 21861
rect 12366 21861 12367 22039
rect 12545 21861 12546 22039
rect 16366 22039 16546 22040
rect 15734 21984 15740 21990
rect 15780 21984 15786 21990
rect 15728 21978 15734 21984
rect 15786 21978 15792 21984
rect 15728 21928 15734 21934
rect 15786 21928 15792 21934
rect 15734 21922 15740 21928
rect 15780 21922 15786 21928
rect 12366 21860 12546 21861
rect 16366 21861 16367 22039
rect 16545 21861 16546 22039
rect 20366 22039 20546 22040
rect 19734 21984 19740 21990
rect 19780 21984 19786 21990
rect 19728 21978 19734 21984
rect 19786 21978 19792 21984
rect 19728 21928 19734 21934
rect 19786 21928 19792 21934
rect 19734 21922 19740 21928
rect 19780 21922 19786 21928
rect 16366 21860 16546 21861
rect 20366 21861 20367 22039
rect 20545 21861 20546 22039
rect 24366 22039 24546 22040
rect 23734 21984 23740 21990
rect 23780 21984 23786 21990
rect 23728 21978 23734 21984
rect 23786 21978 23792 21984
rect 23728 21928 23734 21934
rect 23786 21928 23792 21934
rect 23734 21922 23740 21928
rect 23780 21922 23786 21928
rect 20366 21860 20546 21861
rect 24366 21861 24367 22039
rect 24545 21861 24546 22039
rect 28366 22039 28546 22040
rect 27734 21984 27740 21990
rect 27780 21984 27786 21990
rect 27728 21978 27734 21984
rect 27786 21978 27792 21984
rect 27728 21928 27734 21934
rect 27786 21928 27792 21934
rect 27734 21922 27740 21928
rect 27780 21922 27786 21928
rect 24366 21860 24546 21861
rect 28366 21861 28367 22039
rect 28545 21861 28546 22039
rect 32366 22039 32546 22040
rect 31734 21984 31740 21990
rect 31780 21984 31786 21990
rect 31728 21978 31734 21984
rect 31786 21978 31792 21984
rect 31728 21928 31734 21934
rect 31786 21928 31792 21934
rect 31734 21922 31740 21928
rect 31780 21922 31786 21928
rect 28366 21860 28546 21861
rect 32366 21861 32367 22039
rect 32545 21861 32546 22039
rect 36366 22039 36546 22040
rect 35734 21984 35740 21990
rect 35780 21984 35786 21990
rect 35728 21978 35734 21984
rect 35786 21978 35792 21984
rect 35728 21928 35734 21934
rect 35786 21928 35792 21934
rect 35734 21922 35740 21928
rect 35780 21922 35786 21928
rect 32366 21860 32546 21861
rect 36366 21861 36367 22039
rect 36545 21861 36546 22039
rect 39734 21984 39740 21990
rect 39780 21984 39786 21990
rect 39728 21978 39734 21984
rect 39786 21978 39792 21984
rect 39728 21928 39734 21934
rect 39786 21928 39792 21934
rect 39734 21922 39740 21928
rect 39780 21922 39786 21928
rect 36366 21860 36546 21861
rect 3262 21808 3268 21814
rect 3308 21808 3314 21814
rect 7262 21808 7268 21814
rect 7308 21808 7314 21814
rect 11262 21808 11268 21814
rect 11308 21808 11314 21814
rect 15262 21808 15268 21814
rect 15308 21808 15314 21814
rect 19262 21808 19268 21814
rect 19308 21808 19314 21814
rect 23262 21808 23268 21814
rect 23308 21808 23314 21814
rect 27262 21808 27268 21814
rect 27308 21808 27314 21814
rect 31262 21808 31268 21814
rect 31308 21808 31314 21814
rect 35262 21808 35268 21814
rect 35308 21808 35314 21814
rect 39262 21808 39268 21814
rect 39308 21808 39314 21814
rect 3256 21802 3262 21808
rect 3314 21802 3320 21808
rect 7256 21802 7262 21808
rect 7314 21802 7320 21808
rect 11256 21802 11262 21808
rect 11314 21802 11320 21808
rect 15256 21802 15262 21808
rect 15314 21802 15320 21808
rect 19256 21802 19262 21808
rect 19314 21802 19320 21808
rect 23256 21802 23262 21808
rect 23314 21802 23320 21808
rect 27256 21802 27262 21808
rect 27314 21802 27320 21808
rect 31256 21802 31262 21808
rect 31314 21802 31320 21808
rect 35256 21802 35262 21808
rect 35314 21802 35320 21808
rect 39256 21802 39262 21808
rect 39314 21802 39320 21808
rect 3256 21756 3262 21762
rect 3314 21756 3320 21762
rect 7256 21756 7262 21762
rect 7314 21756 7320 21762
rect 11256 21756 11262 21762
rect 11314 21756 11320 21762
rect 15256 21756 15262 21762
rect 15314 21756 15320 21762
rect 19256 21756 19262 21762
rect 19314 21756 19320 21762
rect 23256 21756 23262 21762
rect 23314 21756 23320 21762
rect 27256 21756 27262 21762
rect 27314 21756 27320 21762
rect 31256 21756 31262 21762
rect 31314 21756 31320 21762
rect 35256 21756 35262 21762
rect 35314 21756 35320 21762
rect 39256 21756 39262 21762
rect 39314 21756 39320 21762
rect 3262 21750 3268 21756
rect 3308 21750 3314 21756
rect 7262 21750 7268 21756
rect 7308 21750 7314 21756
rect 11262 21750 11268 21756
rect 11308 21750 11314 21756
rect 15262 21750 15268 21756
rect 15308 21750 15314 21756
rect 19262 21750 19268 21756
rect 19308 21750 19314 21756
rect 23262 21750 23268 21756
rect 23308 21750 23314 21756
rect 27262 21750 27268 21756
rect 27308 21750 27314 21756
rect 31262 21750 31268 21756
rect 31308 21750 31314 21756
rect 35262 21750 35268 21756
rect 35308 21750 35314 21756
rect 39262 21750 39268 21756
rect 39308 21750 39314 21756
rect 2386 21296 2626 21320
rect 2386 21104 2410 21296
rect 2602 21104 2626 21296
rect 2386 21080 2626 21104
rect 6386 21296 6626 21320
rect 6386 21104 6410 21296
rect 6602 21104 6626 21296
rect 6386 21080 6626 21104
rect 10386 21296 10626 21320
rect 10386 21104 10410 21296
rect 10602 21104 10626 21296
rect 10386 21080 10626 21104
rect 14386 21296 14626 21320
rect 14386 21104 14410 21296
rect 14602 21104 14626 21296
rect 14386 21080 14626 21104
rect 18386 21296 18626 21320
rect 18386 21104 18410 21296
rect 18602 21104 18626 21296
rect 18386 21080 18626 21104
rect 22386 21296 22626 21320
rect 22386 21104 22410 21296
rect 22602 21104 22626 21296
rect 22386 21080 22626 21104
rect 26386 21296 26626 21320
rect 26386 21104 26410 21296
rect 26602 21104 26626 21296
rect 26386 21080 26626 21104
rect 30386 21296 30626 21320
rect 30386 21104 30410 21296
rect 30602 21104 30626 21296
rect 30386 21080 30626 21104
rect 34386 21296 34626 21320
rect 34386 21104 34410 21296
rect 34602 21104 34626 21296
rect 34386 21080 34626 21104
rect 38386 21296 38626 21320
rect 38386 21104 38410 21296
rect 38602 21104 38626 21296
rect 38386 21080 38626 21104
rect 1982 20160 2302 20230
rect 366 19916 606 19940
rect 366 19724 390 19916
rect 582 19724 606 19916
rect 1982 19920 2006 20160
rect 2232 19920 2246 20160
rect 2256 19920 2302 20160
rect 5982 20160 6302 20230
rect 1982 19896 2302 19920
rect 4366 19916 4606 19940
rect 366 19700 606 19724
rect 4366 19724 4390 19916
rect 4582 19724 4606 19916
rect 5982 19920 6006 20160
rect 6232 19920 6246 20160
rect 6256 19920 6302 20160
rect 9982 20160 10302 20230
rect 5982 19896 6302 19920
rect 8366 19916 8606 19940
rect 2852 19709 2996 19714
rect 2852 19639 2857 19709
rect 2991 19639 2996 19709
rect 4366 19700 4606 19724
rect 8366 19724 8390 19916
rect 8582 19724 8606 19916
rect 9982 19920 10006 20160
rect 10232 19920 10246 20160
rect 10256 19920 10302 20160
rect 13982 20160 14302 20230
rect 9982 19896 10302 19920
rect 12366 19916 12606 19940
rect 6852 19709 6996 19714
rect 2852 19634 2996 19639
rect 6852 19639 6857 19709
rect 6991 19639 6996 19709
rect 8366 19700 8606 19724
rect 12366 19724 12390 19916
rect 12582 19724 12606 19916
rect 13982 19920 14006 20160
rect 14232 19920 14246 20160
rect 14256 19920 14302 20160
rect 17982 20160 18302 20230
rect 13982 19896 14302 19920
rect 16366 19916 16606 19940
rect 10852 19709 10996 19714
rect 6852 19634 6996 19639
rect 10852 19639 10857 19709
rect 10991 19639 10996 19709
rect 12366 19700 12606 19724
rect 16366 19724 16390 19916
rect 16582 19724 16606 19916
rect 17982 19920 18006 20160
rect 18232 19920 18246 20160
rect 18256 19920 18302 20160
rect 21982 20160 22302 20230
rect 17982 19896 18302 19920
rect 20366 19916 20606 19940
rect 14852 19709 14996 19714
rect 10852 19634 10996 19639
rect 14852 19639 14857 19709
rect 14991 19639 14996 19709
rect 16366 19700 16606 19724
rect 20366 19724 20390 19916
rect 20582 19724 20606 19916
rect 21982 19920 22006 20160
rect 22232 19920 22246 20160
rect 22256 19920 22302 20160
rect 25982 20160 26302 20230
rect 21982 19896 22302 19920
rect 24366 19916 24606 19940
rect 18852 19709 18996 19714
rect 14852 19634 14996 19639
rect 18852 19639 18857 19709
rect 18991 19639 18996 19709
rect 20366 19700 20606 19724
rect 24366 19724 24390 19916
rect 24582 19724 24606 19916
rect 25982 19920 26006 20160
rect 26232 19920 26246 20160
rect 26256 19920 26302 20160
rect 29982 20160 30302 20230
rect 25982 19896 26302 19920
rect 28366 19916 28606 19940
rect 22852 19709 22996 19714
rect 18852 19634 18996 19639
rect 22852 19639 22857 19709
rect 22991 19639 22996 19709
rect 24366 19700 24606 19724
rect 28366 19724 28390 19916
rect 28582 19724 28606 19916
rect 29982 19920 30006 20160
rect 30232 19920 30246 20160
rect 30256 19920 30302 20160
rect 33982 20160 34302 20230
rect 29982 19896 30302 19920
rect 32366 19916 32606 19940
rect 26852 19709 26996 19714
rect 22852 19634 22996 19639
rect 26852 19639 26857 19709
rect 26991 19639 26996 19709
rect 28366 19700 28606 19724
rect 32366 19724 32390 19916
rect 32582 19724 32606 19916
rect 33982 19920 34006 20160
rect 34232 19920 34246 20160
rect 34256 19920 34302 20160
rect 37982 20160 38302 20230
rect 33982 19896 34302 19920
rect 36366 19916 36606 19940
rect 30852 19709 30996 19714
rect 26852 19634 26996 19639
rect 30852 19639 30857 19709
rect 30991 19639 30996 19709
rect 32366 19700 32606 19724
rect 36366 19724 36390 19916
rect 36582 19724 36606 19916
rect 37982 19920 38006 20160
rect 38232 19920 38246 20160
rect 38256 19920 38302 20160
rect 37982 19896 38302 19920
rect 34852 19709 34996 19714
rect 30852 19634 30996 19639
rect 34852 19639 34857 19709
rect 34991 19639 34996 19709
rect 36366 19700 36606 19724
rect 38852 19709 38996 19714
rect 34852 19634 34996 19639
rect 38852 19639 38857 19709
rect 38991 19639 38996 19709
rect 38852 19634 38996 19639
rect 2366 19559 2546 19560
rect 2366 19381 2367 19559
rect 2545 19381 2546 19559
rect 2366 19380 2546 19381
rect 6366 19559 6546 19560
rect 6366 19381 6367 19559
rect 6545 19381 6546 19559
rect 6366 19380 6546 19381
rect 10366 19559 10546 19560
rect 10366 19381 10367 19559
rect 10545 19381 10546 19559
rect 10366 19380 10546 19381
rect 14366 19559 14546 19560
rect 14366 19381 14367 19559
rect 14545 19381 14546 19559
rect 14366 19380 14546 19381
rect 18366 19559 18546 19560
rect 18366 19381 18367 19559
rect 18545 19381 18546 19559
rect 18366 19380 18546 19381
rect 22366 19559 22546 19560
rect 22366 19381 22367 19559
rect 22545 19381 22546 19559
rect 22366 19380 22546 19381
rect 26366 19559 26546 19560
rect 26366 19381 26367 19559
rect 26545 19381 26546 19559
rect 26366 19380 26546 19381
rect 30366 19559 30546 19560
rect 30366 19381 30367 19559
rect 30545 19381 30546 19559
rect 30366 19380 30546 19381
rect 34366 19559 34546 19560
rect 34366 19381 34367 19559
rect 34545 19381 34546 19559
rect 34366 19380 34546 19381
rect 38366 19559 38546 19560
rect 38366 19381 38367 19559
rect 38545 19381 38546 19559
rect 38366 19380 38546 19381
rect 366 19039 546 19040
rect 366 18861 367 19039
rect 545 18861 546 19039
rect 4366 19039 4546 19040
rect 3734 18984 3740 18990
rect 3780 18984 3786 18990
rect 3728 18978 3734 18984
rect 3786 18978 3792 18984
rect 3728 18928 3734 18934
rect 3786 18928 3792 18934
rect 3734 18922 3740 18928
rect 3780 18922 3786 18928
rect 366 18860 546 18861
rect 4366 18861 4367 19039
rect 4545 18861 4546 19039
rect 8366 19039 8546 19040
rect 7734 18984 7740 18990
rect 7780 18984 7786 18990
rect 7728 18978 7734 18984
rect 7786 18978 7792 18984
rect 7728 18928 7734 18934
rect 7786 18928 7792 18934
rect 7734 18922 7740 18928
rect 7780 18922 7786 18928
rect 4366 18860 4546 18861
rect 8366 18861 8367 19039
rect 8545 18861 8546 19039
rect 12366 19039 12546 19040
rect 11734 18984 11740 18990
rect 11780 18984 11786 18990
rect 11728 18978 11734 18984
rect 11786 18978 11792 18984
rect 11728 18928 11734 18934
rect 11786 18928 11792 18934
rect 11734 18922 11740 18928
rect 11780 18922 11786 18928
rect 8366 18860 8546 18861
rect 12366 18861 12367 19039
rect 12545 18861 12546 19039
rect 16366 19039 16546 19040
rect 15734 18984 15740 18990
rect 15780 18984 15786 18990
rect 15728 18978 15734 18984
rect 15786 18978 15792 18984
rect 15728 18928 15734 18934
rect 15786 18928 15792 18934
rect 15734 18922 15740 18928
rect 15780 18922 15786 18928
rect 12366 18860 12546 18861
rect 16366 18861 16367 19039
rect 16545 18861 16546 19039
rect 20366 19039 20546 19040
rect 19734 18984 19740 18990
rect 19780 18984 19786 18990
rect 19728 18978 19734 18984
rect 19786 18978 19792 18984
rect 19728 18928 19734 18934
rect 19786 18928 19792 18934
rect 19734 18922 19740 18928
rect 19780 18922 19786 18928
rect 16366 18860 16546 18861
rect 20366 18861 20367 19039
rect 20545 18861 20546 19039
rect 24366 19039 24546 19040
rect 23734 18984 23740 18990
rect 23780 18984 23786 18990
rect 23728 18978 23734 18984
rect 23786 18978 23792 18984
rect 23728 18928 23734 18934
rect 23786 18928 23792 18934
rect 23734 18922 23740 18928
rect 23780 18922 23786 18928
rect 20366 18860 20546 18861
rect 24366 18861 24367 19039
rect 24545 18861 24546 19039
rect 28366 19039 28546 19040
rect 27734 18984 27740 18990
rect 27780 18984 27786 18990
rect 27728 18978 27734 18984
rect 27786 18978 27792 18984
rect 27728 18928 27734 18934
rect 27786 18928 27792 18934
rect 27734 18922 27740 18928
rect 27780 18922 27786 18928
rect 24366 18860 24546 18861
rect 28366 18861 28367 19039
rect 28545 18861 28546 19039
rect 32366 19039 32546 19040
rect 31734 18984 31740 18990
rect 31780 18984 31786 18990
rect 31728 18978 31734 18984
rect 31786 18978 31792 18984
rect 31728 18928 31734 18934
rect 31786 18928 31792 18934
rect 31734 18922 31740 18928
rect 31780 18922 31786 18928
rect 28366 18860 28546 18861
rect 32366 18861 32367 19039
rect 32545 18861 32546 19039
rect 36366 19039 36546 19040
rect 35734 18984 35740 18990
rect 35780 18984 35786 18990
rect 35728 18978 35734 18984
rect 35786 18978 35792 18984
rect 35728 18928 35734 18934
rect 35786 18928 35792 18934
rect 35734 18922 35740 18928
rect 35780 18922 35786 18928
rect 32366 18860 32546 18861
rect 36366 18861 36367 19039
rect 36545 18861 36546 19039
rect 39734 18984 39740 18990
rect 39780 18984 39786 18990
rect 39728 18978 39734 18984
rect 39786 18978 39792 18984
rect 39728 18928 39734 18934
rect 39786 18928 39792 18934
rect 39734 18922 39740 18928
rect 39780 18922 39786 18928
rect 36366 18860 36546 18861
rect 3262 18808 3268 18814
rect 3308 18808 3314 18814
rect 7262 18808 7268 18814
rect 7308 18808 7314 18814
rect 11262 18808 11268 18814
rect 11308 18808 11314 18814
rect 15262 18808 15268 18814
rect 15308 18808 15314 18814
rect 19262 18808 19268 18814
rect 19308 18808 19314 18814
rect 23262 18808 23268 18814
rect 23308 18808 23314 18814
rect 27262 18808 27268 18814
rect 27308 18808 27314 18814
rect 31262 18808 31268 18814
rect 31308 18808 31314 18814
rect 35262 18808 35268 18814
rect 35308 18808 35314 18814
rect 39262 18808 39268 18814
rect 39308 18808 39314 18814
rect 3256 18802 3262 18808
rect 3314 18802 3320 18808
rect 7256 18802 7262 18808
rect 7314 18802 7320 18808
rect 11256 18802 11262 18808
rect 11314 18802 11320 18808
rect 15256 18802 15262 18808
rect 15314 18802 15320 18808
rect 19256 18802 19262 18808
rect 19314 18802 19320 18808
rect 23256 18802 23262 18808
rect 23314 18802 23320 18808
rect 27256 18802 27262 18808
rect 27314 18802 27320 18808
rect 31256 18802 31262 18808
rect 31314 18802 31320 18808
rect 35256 18802 35262 18808
rect 35314 18802 35320 18808
rect 39256 18802 39262 18808
rect 39314 18802 39320 18808
rect 3256 18756 3262 18762
rect 3314 18756 3320 18762
rect 7256 18756 7262 18762
rect 7314 18756 7320 18762
rect 11256 18756 11262 18762
rect 11314 18756 11320 18762
rect 15256 18756 15262 18762
rect 15314 18756 15320 18762
rect 19256 18756 19262 18762
rect 19314 18756 19320 18762
rect 23256 18756 23262 18762
rect 23314 18756 23320 18762
rect 27256 18756 27262 18762
rect 27314 18756 27320 18762
rect 31256 18756 31262 18762
rect 31314 18756 31320 18762
rect 35256 18756 35262 18762
rect 35314 18756 35320 18762
rect 39256 18756 39262 18762
rect 39314 18756 39320 18762
rect 3262 18750 3268 18756
rect 3308 18750 3314 18756
rect 7262 18750 7268 18756
rect 7308 18750 7314 18756
rect 11262 18750 11268 18756
rect 11308 18750 11314 18756
rect 15262 18750 15268 18756
rect 15308 18750 15314 18756
rect 19262 18750 19268 18756
rect 19308 18750 19314 18756
rect 23262 18750 23268 18756
rect 23308 18750 23314 18756
rect 27262 18750 27268 18756
rect 27308 18750 27314 18756
rect 31262 18750 31268 18756
rect 31308 18750 31314 18756
rect 35262 18750 35268 18756
rect 35308 18750 35314 18756
rect 39262 18750 39268 18756
rect 39308 18750 39314 18756
rect 2386 18296 2626 18320
rect 2386 18104 2410 18296
rect 2602 18104 2626 18296
rect 2386 18080 2626 18104
rect 6386 18296 6626 18320
rect 6386 18104 6410 18296
rect 6602 18104 6626 18296
rect 6386 18080 6626 18104
rect 10386 18296 10626 18320
rect 10386 18104 10410 18296
rect 10602 18104 10626 18296
rect 10386 18080 10626 18104
rect 14386 18296 14626 18320
rect 14386 18104 14410 18296
rect 14602 18104 14626 18296
rect 14386 18080 14626 18104
rect 18386 18296 18626 18320
rect 18386 18104 18410 18296
rect 18602 18104 18626 18296
rect 18386 18080 18626 18104
rect 22386 18296 22626 18320
rect 22386 18104 22410 18296
rect 22602 18104 22626 18296
rect 22386 18080 22626 18104
rect 26386 18296 26626 18320
rect 26386 18104 26410 18296
rect 26602 18104 26626 18296
rect 26386 18080 26626 18104
rect 30386 18296 30626 18320
rect 30386 18104 30410 18296
rect 30602 18104 30626 18296
rect 30386 18080 30626 18104
rect 34386 18296 34626 18320
rect 34386 18104 34410 18296
rect 34602 18104 34626 18296
rect 34386 18080 34626 18104
rect 38386 18296 38626 18320
rect 38386 18104 38410 18296
rect 38602 18104 38626 18296
rect 38386 18080 38626 18104
rect 1982 17160 2302 17230
rect 366 16916 606 16940
rect 366 16724 390 16916
rect 582 16724 606 16916
rect 1982 16920 2006 17160
rect 2232 16920 2246 17160
rect 2256 16920 2302 17160
rect 5982 17160 6302 17230
rect 1982 16896 2302 16920
rect 4366 16916 4606 16940
rect 366 16700 606 16724
rect 4366 16724 4390 16916
rect 4582 16724 4606 16916
rect 5982 16920 6006 17160
rect 6232 16920 6246 17160
rect 6256 16920 6302 17160
rect 9982 17160 10302 17230
rect 5982 16896 6302 16920
rect 8366 16916 8606 16940
rect 2852 16709 2996 16714
rect 2852 16639 2857 16709
rect 2991 16639 2996 16709
rect 4366 16700 4606 16724
rect 8366 16724 8390 16916
rect 8582 16724 8606 16916
rect 9982 16920 10006 17160
rect 10232 16920 10246 17160
rect 10256 16920 10302 17160
rect 13982 17160 14302 17230
rect 9982 16896 10302 16920
rect 12366 16916 12606 16940
rect 6852 16709 6996 16714
rect 2852 16634 2996 16639
rect 6852 16639 6857 16709
rect 6991 16639 6996 16709
rect 8366 16700 8606 16724
rect 12366 16724 12390 16916
rect 12582 16724 12606 16916
rect 13982 16920 14006 17160
rect 14232 16920 14246 17160
rect 14256 16920 14302 17160
rect 17982 17160 18302 17230
rect 13982 16896 14302 16920
rect 16366 16916 16606 16940
rect 10852 16709 10996 16714
rect 6852 16634 6996 16639
rect 10852 16639 10857 16709
rect 10991 16639 10996 16709
rect 12366 16700 12606 16724
rect 16366 16724 16390 16916
rect 16582 16724 16606 16916
rect 17982 16920 18006 17160
rect 18232 16920 18246 17160
rect 18256 16920 18302 17160
rect 21982 17160 22302 17230
rect 17982 16896 18302 16920
rect 20366 16916 20606 16940
rect 14852 16709 14996 16714
rect 10852 16634 10996 16639
rect 14852 16639 14857 16709
rect 14991 16639 14996 16709
rect 16366 16700 16606 16724
rect 20366 16724 20390 16916
rect 20582 16724 20606 16916
rect 21982 16920 22006 17160
rect 22232 16920 22246 17160
rect 22256 16920 22302 17160
rect 25982 17160 26302 17230
rect 21982 16896 22302 16920
rect 24366 16916 24606 16940
rect 18852 16709 18996 16714
rect 14852 16634 14996 16639
rect 18852 16639 18857 16709
rect 18991 16639 18996 16709
rect 20366 16700 20606 16724
rect 24366 16724 24390 16916
rect 24582 16724 24606 16916
rect 25982 16920 26006 17160
rect 26232 16920 26246 17160
rect 26256 16920 26302 17160
rect 29982 17160 30302 17230
rect 25982 16896 26302 16920
rect 28366 16916 28606 16940
rect 22852 16709 22996 16714
rect 18852 16634 18996 16639
rect 22852 16639 22857 16709
rect 22991 16639 22996 16709
rect 24366 16700 24606 16724
rect 28366 16724 28390 16916
rect 28582 16724 28606 16916
rect 29982 16920 30006 17160
rect 30232 16920 30246 17160
rect 30256 16920 30302 17160
rect 33982 17160 34302 17230
rect 29982 16896 30302 16920
rect 32366 16916 32606 16940
rect 26852 16709 26996 16714
rect 22852 16634 22996 16639
rect 26852 16639 26857 16709
rect 26991 16639 26996 16709
rect 28366 16700 28606 16724
rect 32366 16724 32390 16916
rect 32582 16724 32606 16916
rect 33982 16920 34006 17160
rect 34232 16920 34246 17160
rect 34256 16920 34302 17160
rect 37982 17160 38302 17230
rect 33982 16896 34302 16920
rect 36366 16916 36606 16940
rect 30852 16709 30996 16714
rect 26852 16634 26996 16639
rect 30852 16639 30857 16709
rect 30991 16639 30996 16709
rect 32366 16700 32606 16724
rect 36366 16724 36390 16916
rect 36582 16724 36606 16916
rect 37982 16920 38006 17160
rect 38232 16920 38246 17160
rect 38256 16920 38302 17160
rect 37982 16896 38302 16920
rect 34852 16709 34996 16714
rect 30852 16634 30996 16639
rect 34852 16639 34857 16709
rect 34991 16639 34996 16709
rect 36366 16700 36606 16724
rect 38852 16709 38996 16714
rect 34852 16634 34996 16639
rect 38852 16639 38857 16709
rect 38991 16639 38996 16709
rect 38852 16634 38996 16639
rect 2366 16559 2546 16560
rect 2366 16381 2367 16559
rect 2545 16381 2546 16559
rect 2366 16380 2546 16381
rect 6366 16559 6546 16560
rect 6366 16381 6367 16559
rect 6545 16381 6546 16559
rect 6366 16380 6546 16381
rect 10366 16559 10546 16560
rect 10366 16381 10367 16559
rect 10545 16381 10546 16559
rect 10366 16380 10546 16381
rect 14366 16559 14546 16560
rect 14366 16381 14367 16559
rect 14545 16381 14546 16559
rect 14366 16380 14546 16381
rect 18366 16559 18546 16560
rect 18366 16381 18367 16559
rect 18545 16381 18546 16559
rect 18366 16380 18546 16381
rect 22366 16559 22546 16560
rect 22366 16381 22367 16559
rect 22545 16381 22546 16559
rect 22366 16380 22546 16381
rect 26366 16559 26546 16560
rect 26366 16381 26367 16559
rect 26545 16381 26546 16559
rect 26366 16380 26546 16381
rect 30366 16559 30546 16560
rect 30366 16381 30367 16559
rect 30545 16381 30546 16559
rect 30366 16380 30546 16381
rect 34366 16559 34546 16560
rect 34366 16381 34367 16559
rect 34545 16381 34546 16559
rect 34366 16380 34546 16381
rect 38366 16559 38546 16560
rect 38366 16381 38367 16559
rect 38545 16381 38546 16559
rect 38366 16380 38546 16381
rect 366 16039 546 16040
rect 366 15861 367 16039
rect 545 15861 546 16039
rect 4366 16039 4546 16040
rect 3734 15984 3740 15990
rect 3780 15984 3786 15990
rect 3728 15978 3734 15984
rect 3786 15978 3792 15984
rect 3728 15928 3734 15934
rect 3786 15928 3792 15934
rect 3734 15922 3740 15928
rect 3780 15922 3786 15928
rect 366 15860 546 15861
rect 4366 15861 4367 16039
rect 4545 15861 4546 16039
rect 8366 16039 8546 16040
rect 7734 15984 7740 15990
rect 7780 15984 7786 15990
rect 7728 15978 7734 15984
rect 7786 15978 7792 15984
rect 7728 15928 7734 15934
rect 7786 15928 7792 15934
rect 7734 15922 7740 15928
rect 7780 15922 7786 15928
rect 4366 15860 4546 15861
rect 8366 15861 8367 16039
rect 8545 15861 8546 16039
rect 12366 16039 12546 16040
rect 11734 15984 11740 15990
rect 11780 15984 11786 15990
rect 11728 15978 11734 15984
rect 11786 15978 11792 15984
rect 11728 15928 11734 15934
rect 11786 15928 11792 15934
rect 11734 15922 11740 15928
rect 11780 15922 11786 15928
rect 8366 15860 8546 15861
rect 12366 15861 12367 16039
rect 12545 15861 12546 16039
rect 16366 16039 16546 16040
rect 15734 15984 15740 15990
rect 15780 15984 15786 15990
rect 15728 15978 15734 15984
rect 15786 15978 15792 15984
rect 15728 15928 15734 15934
rect 15786 15928 15792 15934
rect 15734 15922 15740 15928
rect 15780 15922 15786 15928
rect 12366 15860 12546 15861
rect 16366 15861 16367 16039
rect 16545 15861 16546 16039
rect 20366 16039 20546 16040
rect 19734 15984 19740 15990
rect 19780 15984 19786 15990
rect 19728 15978 19734 15984
rect 19786 15978 19792 15984
rect 19728 15928 19734 15934
rect 19786 15928 19792 15934
rect 19734 15922 19740 15928
rect 19780 15922 19786 15928
rect 16366 15860 16546 15861
rect 20366 15861 20367 16039
rect 20545 15861 20546 16039
rect 24366 16039 24546 16040
rect 23734 15984 23740 15990
rect 23780 15984 23786 15990
rect 23728 15978 23734 15984
rect 23786 15978 23792 15984
rect 23728 15928 23734 15934
rect 23786 15928 23792 15934
rect 23734 15922 23740 15928
rect 23780 15922 23786 15928
rect 20366 15860 20546 15861
rect 24366 15861 24367 16039
rect 24545 15861 24546 16039
rect 28366 16039 28546 16040
rect 27734 15984 27740 15990
rect 27780 15984 27786 15990
rect 27728 15978 27734 15984
rect 27786 15978 27792 15984
rect 27728 15928 27734 15934
rect 27786 15928 27792 15934
rect 27734 15922 27740 15928
rect 27780 15922 27786 15928
rect 24366 15860 24546 15861
rect 28366 15861 28367 16039
rect 28545 15861 28546 16039
rect 32366 16039 32546 16040
rect 31734 15984 31740 15990
rect 31780 15984 31786 15990
rect 31728 15978 31734 15984
rect 31786 15978 31792 15984
rect 31728 15928 31734 15934
rect 31786 15928 31792 15934
rect 31734 15922 31740 15928
rect 31780 15922 31786 15928
rect 28366 15860 28546 15861
rect 32366 15861 32367 16039
rect 32545 15861 32546 16039
rect 36366 16039 36546 16040
rect 35734 15984 35740 15990
rect 35780 15984 35786 15990
rect 35728 15978 35734 15984
rect 35786 15978 35792 15984
rect 35728 15928 35734 15934
rect 35786 15928 35792 15934
rect 35734 15922 35740 15928
rect 35780 15922 35786 15928
rect 32366 15860 32546 15861
rect 36366 15861 36367 16039
rect 36545 15861 36546 16039
rect 39734 15984 39740 15990
rect 39780 15984 39786 15990
rect 39728 15978 39734 15984
rect 39786 15978 39792 15984
rect 39728 15928 39734 15934
rect 39786 15928 39792 15934
rect 39734 15922 39740 15928
rect 39780 15922 39786 15928
rect 36366 15860 36546 15861
rect 3262 15808 3268 15814
rect 3308 15808 3314 15814
rect 7262 15808 7268 15814
rect 7308 15808 7314 15814
rect 11262 15808 11268 15814
rect 11308 15808 11314 15814
rect 15262 15808 15268 15814
rect 15308 15808 15314 15814
rect 19262 15808 19268 15814
rect 19308 15808 19314 15814
rect 23262 15808 23268 15814
rect 23308 15808 23314 15814
rect 27262 15808 27268 15814
rect 27308 15808 27314 15814
rect 31262 15808 31268 15814
rect 31308 15808 31314 15814
rect 35262 15808 35268 15814
rect 35308 15808 35314 15814
rect 39262 15808 39268 15814
rect 39308 15808 39314 15814
rect 3256 15802 3262 15808
rect 3314 15802 3320 15808
rect 7256 15802 7262 15808
rect 7314 15802 7320 15808
rect 11256 15802 11262 15808
rect 11314 15802 11320 15808
rect 15256 15802 15262 15808
rect 15314 15802 15320 15808
rect 19256 15802 19262 15808
rect 19314 15802 19320 15808
rect 23256 15802 23262 15808
rect 23314 15802 23320 15808
rect 27256 15802 27262 15808
rect 27314 15802 27320 15808
rect 31256 15802 31262 15808
rect 31314 15802 31320 15808
rect 35256 15802 35262 15808
rect 35314 15802 35320 15808
rect 39256 15802 39262 15808
rect 39314 15802 39320 15808
rect 3256 15756 3262 15762
rect 3314 15756 3320 15762
rect 7256 15756 7262 15762
rect 7314 15756 7320 15762
rect 11256 15756 11262 15762
rect 11314 15756 11320 15762
rect 15256 15756 15262 15762
rect 15314 15756 15320 15762
rect 19256 15756 19262 15762
rect 19314 15756 19320 15762
rect 23256 15756 23262 15762
rect 23314 15756 23320 15762
rect 27256 15756 27262 15762
rect 27314 15756 27320 15762
rect 31256 15756 31262 15762
rect 31314 15756 31320 15762
rect 35256 15756 35262 15762
rect 35314 15756 35320 15762
rect 39256 15756 39262 15762
rect 39314 15756 39320 15762
rect 3262 15750 3268 15756
rect 3308 15750 3314 15756
rect 7262 15750 7268 15756
rect 7308 15750 7314 15756
rect 11262 15750 11268 15756
rect 11308 15750 11314 15756
rect 15262 15750 15268 15756
rect 15308 15750 15314 15756
rect 19262 15750 19268 15756
rect 19308 15750 19314 15756
rect 23262 15750 23268 15756
rect 23308 15750 23314 15756
rect 27262 15750 27268 15756
rect 27308 15750 27314 15756
rect 31262 15750 31268 15756
rect 31308 15750 31314 15756
rect 35262 15750 35268 15756
rect 35308 15750 35314 15756
rect 39262 15750 39268 15756
rect 39308 15750 39314 15756
rect 4366 13724 4390 13740
rect 4582 13724 4606 13740
rect 2856 13711 2992 13716
rect 2856 13637 2861 13711
rect 2987 13637 2992 13711
rect 4366 13700 4606 13724
rect 38856 13711 38992 13716
rect 2856 13632 2992 13637
rect 38856 13637 38861 13711
rect 38987 13637 38992 13711
rect 38856 13632 38992 13637
rect 2366 13559 2546 13560
rect 2366 13381 2367 13559
rect 2545 13381 2546 13559
rect 2366 13380 2546 13381
rect 6366 13559 6486 13560
rect 38366 13559 38546 13560
rect 6366 13381 6367 13559
rect 38366 13381 38367 13559
rect 38545 13381 38546 13559
rect 6366 13380 6486 13381
rect 38366 13380 38546 13381
rect 3728 13010 3734 13016
rect 3780 13010 3786 13016
rect 39728 13010 39734 13016
rect 39780 13010 39786 13016
rect 3722 13004 3728 13010
rect 3786 13004 3792 13010
rect 39722 13004 39728 13010
rect 39786 13004 39792 13010
rect 4386 12999 4566 13000
rect 3722 12948 3728 12954
rect 3786 12948 3792 12954
rect 3728 12942 3734 12948
rect 3780 12942 3786 12948
rect 4386 12821 4387 12999
rect 4565 12821 4566 12999
rect 39722 12948 39728 12954
rect 39786 12948 39792 12954
rect 39728 12942 39734 12948
rect 39780 12942 39786 12948
rect 4386 12820 4566 12821
rect 3262 12808 3268 12814
rect 3308 12808 3314 12814
rect 39262 12808 39268 12814
rect 39308 12808 39314 12814
rect 3256 12802 3262 12808
rect 3314 12802 3320 12808
rect 39256 12802 39262 12808
rect 39314 12802 39320 12808
rect 3256 12756 3262 12762
rect 3314 12756 3320 12762
rect 39256 12756 39262 12762
rect 39314 12756 39320 12762
rect 3262 12750 3268 12756
rect 3308 12750 3314 12756
rect 39262 12750 39268 12756
rect 39308 12750 39314 12756
rect 2286 12296 2526 12320
rect 2286 12104 2310 12296
rect 2502 12104 2526 12296
rect 2286 12080 2526 12104
rect 6286 12296 6486 12320
rect 38286 12296 38526 12320
rect 6286 12104 6310 12296
rect 38286 12104 38310 12296
rect 38502 12104 38526 12296
rect 6286 12080 6486 12104
rect 38286 12080 38526 12104
rect 1982 11160 2302 11222
rect 1982 10920 2006 11160
rect 2242 10920 2246 11160
rect 2266 10920 2302 11160
rect 5982 11160 6302 11222
rect 1982 10896 2302 10920
rect 4366 10916 4606 10940
rect 4366 10724 4390 10916
rect 4582 10724 4606 10916
rect 5982 10920 6006 11160
rect 6242 10920 6246 11160
rect 6266 10920 6302 11160
rect 5982 10896 6302 10920
rect 37982 11160 38302 11222
rect 37982 10920 38006 11160
rect 38242 10920 38246 11160
rect 38266 10920 38302 11160
rect 37982 10896 38302 10920
rect 2856 10711 2992 10716
rect 2856 10637 2861 10711
rect 2987 10637 2992 10711
rect 4366 10700 4606 10724
rect 38856 10711 38992 10716
rect 2856 10632 2992 10637
rect 38856 10637 38861 10711
rect 38987 10637 38992 10711
rect 38856 10632 38992 10637
rect 2366 10559 2546 10560
rect 2366 10381 2367 10559
rect 2545 10381 2546 10559
rect 2366 10380 2546 10381
rect 6366 10559 6486 10560
rect 38366 10559 38546 10560
rect 6366 10381 6367 10559
rect 38366 10381 38367 10559
rect 38545 10381 38546 10559
rect 6366 10380 6486 10381
rect 38366 10380 38546 10381
rect 3728 10010 3734 10016
rect 3780 10010 3786 10016
rect 39728 10010 39734 10016
rect 39780 10010 39786 10016
rect 3722 10004 3728 10010
rect 3786 10004 3792 10010
rect 39722 10004 39728 10010
rect 39786 10004 39792 10010
rect 4386 9999 4566 10000
rect 3722 9948 3728 9954
rect 3786 9948 3792 9954
rect 3728 9942 3734 9948
rect 3780 9942 3786 9948
rect 4386 9821 4387 9999
rect 4565 9821 4566 9999
rect 39722 9948 39728 9954
rect 39786 9948 39792 9954
rect 39728 9942 39734 9948
rect 39780 9942 39786 9948
rect 4386 9820 4566 9821
rect 3262 9808 3268 9814
rect 3308 9808 3314 9814
rect 39262 9808 39268 9814
rect 39308 9808 39314 9814
rect 3256 9802 3262 9808
rect 3314 9802 3320 9808
rect 39256 9802 39262 9808
rect 39314 9802 39320 9808
rect 3256 9756 3262 9762
rect 3314 9756 3320 9762
rect 39256 9756 39262 9762
rect 39314 9756 39320 9762
rect 3262 9750 3268 9756
rect 3308 9750 3314 9756
rect 39262 9750 39268 9756
rect 39308 9750 39314 9756
rect 2286 9296 2526 9320
rect 2286 9104 2310 9296
rect 2502 9104 2526 9296
rect 2286 9080 2526 9104
rect 6286 9296 6486 9320
rect 38286 9296 38526 9320
rect 6286 9104 6310 9296
rect 38286 9104 38310 9296
rect 38502 9104 38526 9296
rect 6286 9080 6486 9104
rect 38286 9080 38526 9104
rect 1982 8160 2302 8222
rect 1982 7920 2006 8160
rect 2242 7920 2246 8160
rect 2266 7920 2302 8160
rect 5982 8160 6302 8222
rect 1982 7896 2302 7920
rect 4366 7916 4606 7940
rect 4366 7724 4390 7916
rect 4582 7724 4606 7916
rect 5982 7920 6006 8160
rect 6242 7920 6246 8160
rect 6266 7920 6302 8160
rect 5982 7896 6302 7920
rect 37982 8160 38302 8222
rect 37982 7920 38006 8160
rect 38242 7920 38246 8160
rect 38266 7920 38302 8160
rect 37982 7896 38302 7920
rect 2856 7711 2992 7716
rect 2856 7637 2861 7711
rect 2987 7637 2992 7711
rect 4366 7700 4606 7724
rect 38856 7711 38992 7716
rect 2856 7632 2992 7637
rect 38856 7637 38861 7711
rect 38987 7637 38992 7711
rect 38856 7632 38992 7637
rect 2366 7559 2546 7560
rect 2366 7381 2367 7559
rect 2545 7381 2546 7559
rect 2366 7380 2546 7381
rect 6366 7559 6486 7560
rect 38366 7559 38546 7560
rect 6366 7381 6367 7559
rect 38366 7381 38367 7559
rect 38545 7381 38546 7559
rect 6366 7380 6486 7381
rect 38366 7380 38546 7381
rect 3728 7010 3734 7016
rect 3780 7010 3786 7016
rect 39728 7010 39734 7016
rect 39780 7010 39786 7016
rect 3722 7004 3728 7010
rect 3786 7004 3792 7010
rect 39722 7004 39728 7010
rect 39786 7004 39792 7010
rect 4386 6999 4566 7000
rect 3722 6948 3728 6954
rect 3786 6948 3792 6954
rect 3728 6942 3734 6948
rect 3780 6942 3786 6948
rect 4386 6821 4387 6999
rect 4565 6821 4566 6999
rect 39722 6948 39728 6954
rect 39786 6948 39792 6954
rect 39728 6942 39734 6948
rect 39780 6942 39786 6948
rect 4386 6820 4566 6821
rect 3262 6808 3268 6814
rect 3308 6808 3314 6814
rect 39262 6808 39268 6814
rect 39308 6808 39314 6814
rect 3256 6802 3262 6808
rect 3314 6802 3320 6808
rect 39256 6802 39262 6808
rect 39314 6802 39320 6808
rect 3256 6756 3262 6762
rect 3314 6756 3320 6762
rect 39256 6756 39262 6762
rect 39314 6756 39320 6762
rect 3262 6750 3268 6756
rect 3308 6750 3314 6756
rect 39262 6750 39268 6756
rect 39308 6750 39314 6756
rect 2286 6296 2526 6320
rect 2286 6104 2310 6296
rect 2502 6104 2526 6296
rect 2286 6080 2526 6104
rect 6286 6296 6486 6320
rect 38286 6296 38526 6320
rect 6286 6104 6310 6296
rect 38286 6104 38310 6296
rect 38502 6104 38526 6296
rect 6286 6080 6486 6104
rect 38286 6080 38526 6104
rect 1982 5160 2302 5222
rect 1982 4920 2006 5160
rect 2242 4920 2246 5160
rect 2266 4920 2302 5160
rect 5982 5160 6302 5222
rect 1982 4896 2302 4920
rect 4366 4916 4606 4940
rect 4366 4724 4390 4916
rect 4582 4724 4606 4916
rect 5982 4920 6006 5160
rect 6242 4920 6246 5160
rect 6266 4920 6302 5160
rect 5982 4896 6302 4920
rect 37982 5160 38302 5222
rect 37982 4920 38006 5160
rect 38242 4920 38246 5160
rect 38266 4920 38302 5160
rect 37982 4896 38302 4920
rect 2856 4711 2992 4716
rect 2856 4637 2861 4711
rect 2987 4637 2992 4711
rect 4366 4700 4606 4724
rect 38856 4711 38992 4716
rect 2856 4632 2992 4637
rect 38856 4637 38861 4711
rect 38987 4637 38992 4711
rect 38856 4632 38992 4637
rect 2366 4559 2546 4560
rect 2366 4381 2367 4559
rect 2545 4381 2546 4559
rect 2366 4380 2546 4381
rect 6366 4559 6486 4560
rect 38366 4559 38546 4560
rect 6366 4381 6367 4559
rect 38366 4381 38367 4559
rect 38545 4381 38546 4559
rect 6366 4380 6486 4381
rect 38366 4380 38546 4381
rect 3728 4010 3734 4016
rect 3780 4010 3786 4016
rect 39728 4010 39734 4016
rect 39780 4010 39786 4016
rect 3722 4004 3728 4010
rect 3786 4004 3792 4010
rect 39722 4004 39728 4010
rect 39786 4004 39792 4010
rect 4386 3999 4566 4000
rect 3722 3948 3728 3954
rect 3786 3948 3792 3954
rect 3728 3942 3734 3948
rect 3780 3942 3786 3948
rect 4386 3821 4387 3999
rect 4565 3821 4566 3999
rect 39722 3948 39728 3954
rect 39786 3948 39792 3954
rect 39728 3942 39734 3948
rect 39780 3942 39786 3948
rect 4386 3820 4566 3821
rect 3262 3808 3268 3814
rect 3308 3808 3314 3814
rect 39262 3808 39268 3814
rect 39308 3808 39314 3814
rect 3256 3802 3262 3808
rect 3314 3802 3320 3808
rect 39256 3802 39262 3808
rect 39314 3802 39320 3808
rect 3256 3756 3262 3762
rect 3314 3756 3320 3762
rect 39256 3756 39262 3762
rect 39314 3756 39320 3762
rect 3262 3750 3268 3756
rect 3308 3750 3314 3756
rect 39262 3750 39268 3756
rect 39308 3750 39314 3756
rect 2286 3296 2526 3320
rect 2286 3104 2310 3296
rect 2502 3104 2526 3296
rect 2286 3080 2526 3104
rect 6286 3296 6486 3320
rect 38286 3296 38526 3320
rect 6286 3104 6310 3296
rect 38286 3104 38310 3296
rect 38502 3104 38526 3296
rect 6286 3080 6486 3104
rect 38286 3080 38526 3104
rect 1982 2160 2302 2222
rect 1982 1920 2006 2160
rect 2242 1920 2246 2160
rect 2266 1920 2302 2160
rect 5982 2160 6302 2222
rect 1982 1896 2302 1920
rect 4366 1916 4606 1940
rect 4366 1724 4390 1916
rect 4582 1724 4606 1916
rect 5982 1920 6006 2160
rect 6242 1920 6246 2160
rect 6266 1920 6302 2160
rect 5982 1896 6302 1920
rect 37982 2160 38302 2222
rect 37982 1920 38006 2160
rect 38242 1920 38246 2160
rect 38266 1920 38302 2160
rect 37982 1896 38302 1920
rect 2856 1711 2992 1716
rect 2856 1637 2861 1711
rect 2987 1637 2992 1711
rect 4366 1700 4606 1724
rect 38856 1711 38992 1716
rect 2856 1632 2992 1637
rect 38856 1637 38861 1711
rect 38987 1637 38992 1711
rect 38856 1632 38992 1637
rect 2366 1559 2546 1560
rect 2366 1381 2367 1559
rect 2545 1381 2546 1559
rect 2366 1380 2546 1381
rect 6366 1559 6486 1560
rect 38366 1559 38546 1560
rect 6366 1381 6367 1559
rect 38366 1381 38367 1559
rect 38545 1381 38546 1559
rect 6366 1380 6486 1381
rect 38366 1380 38546 1381
rect 3728 1010 3734 1016
rect 3780 1010 3786 1016
rect 39728 1010 39734 1016
rect 39780 1010 39786 1016
rect 3722 1004 3728 1010
rect 3786 1004 3792 1010
rect 39722 1004 39728 1010
rect 39786 1004 39792 1010
rect 4386 999 4566 1000
rect 3722 948 3728 954
rect 3786 948 3792 954
rect 3728 942 3734 948
rect 3780 942 3786 948
rect 4386 821 4387 999
rect 4565 821 4566 999
rect 39722 948 39728 954
rect 39786 948 39792 954
rect 39728 942 39734 948
rect 39780 942 39786 948
rect 4386 820 4566 821
rect 3262 808 3268 814
rect 3308 808 3314 814
rect 39262 808 39268 814
rect 39308 808 39314 814
rect 3256 802 3262 808
rect 3314 802 3320 808
rect 39256 802 39262 808
rect 39314 802 39320 808
rect 3256 756 3262 762
rect 3314 756 3320 762
rect 39256 756 39262 762
rect 39314 756 39320 762
rect 3262 750 3268 756
rect 3308 750 3314 756
rect 39262 750 39268 756
rect 39308 750 39314 756
rect 2286 296 2526 320
rect 2286 104 2310 296
rect 2502 104 2526 296
rect 2286 80 2526 104
rect 6286 296 6486 320
rect 38286 296 38526 320
rect 6286 104 6310 296
rect 38286 104 38310 296
rect 38502 104 38526 296
rect 6286 80 6486 104
rect 38286 80 38526 104
<< error_s >>
rect 2386 15296 2626 15320
rect 2386 15104 2410 15296
rect 2602 15104 2626 15296
rect 2386 15080 2626 15104
rect 6386 15296 6626 15320
rect 6386 15104 6410 15296
rect 6602 15104 6626 15296
rect 6386 15080 6626 15104
rect 10386 15296 10626 15320
rect 10386 15104 10410 15296
rect 10602 15104 10626 15296
rect 10386 15080 10626 15104
rect 14386 15296 14626 15320
rect 14386 15104 14410 15296
rect 14602 15104 14626 15296
rect 14386 15080 14626 15104
rect 18386 15296 18626 15320
rect 18386 15104 18410 15296
rect 18602 15104 18626 15296
rect 18386 15080 18626 15104
rect 22386 15296 22626 15320
rect 22386 15104 22410 15296
rect 22602 15104 22626 15296
rect 22386 15080 22626 15104
rect 26386 15296 26626 15320
rect 26386 15104 26410 15296
rect 26602 15104 26626 15296
rect 26386 15080 26626 15104
rect 30386 15296 30626 15320
rect 30386 15104 30410 15296
rect 30602 15104 30626 15296
rect 30386 15080 30626 15104
rect 34386 15296 34626 15320
rect 34386 15104 34410 15296
rect 34602 15104 34626 15296
rect 34386 15080 34626 15104
rect 38386 15296 38626 15320
rect 38386 15104 38410 15296
rect 38602 15104 38626 15296
rect 38386 15080 38626 15104
rect 1982 14160 2302 14222
rect 366 13916 606 13940
rect 366 13740 390 13916
rect 582 13740 606 13916
rect 1982 13920 2006 14160
rect 2242 13920 2246 14160
rect 2266 13920 2302 14160
rect 5982 14160 6302 14222
rect 1982 13896 2302 13920
rect 4366 13916 4606 13940
rect 4366 13740 4390 13916
rect 4582 13740 4606 13916
rect 5982 13920 6006 14160
rect 6242 13920 6246 14160
rect 6266 13920 6302 14160
rect 9982 14160 10302 14222
rect 5982 13896 6302 13920
rect 8366 13916 8606 13940
rect 8366 13740 8390 13916
rect 8582 13740 8606 13916
rect 9982 13920 10006 14160
rect 10242 13920 10246 14160
rect 10266 13920 10302 14160
rect 13982 14160 14302 14222
rect 9982 13896 10302 13920
rect 12366 13916 12606 13940
rect 12366 13740 12390 13916
rect 12582 13740 12606 13916
rect 13982 13920 14006 14160
rect 14242 13920 14246 14160
rect 14266 13920 14302 14160
rect 17982 14160 18302 14222
rect 13982 13896 14302 13920
rect 16366 13916 16606 13940
rect 16366 13740 16390 13916
rect 16582 13740 16606 13916
rect 17982 13920 18006 14160
rect 18242 13920 18246 14160
rect 18266 13920 18302 14160
rect 21982 14160 22302 14222
rect 17982 13896 18302 13920
rect 20366 13916 20606 13940
rect 20366 13740 20390 13916
rect 20582 13740 20606 13916
rect 21982 13920 22006 14160
rect 22242 13920 22246 14160
rect 22266 13920 22302 14160
rect 25982 14160 26302 14222
rect 21982 13896 22302 13920
rect 24366 13916 24606 13940
rect 24366 13740 24390 13916
rect 24582 13740 24606 13916
rect 25982 13920 26006 14160
rect 26242 13920 26246 14160
rect 26266 13920 26302 14160
rect 29982 14160 30302 14222
rect 25982 13896 26302 13920
rect 28366 13916 28606 13940
rect 28366 13740 28390 13916
rect 28582 13740 28606 13916
rect 29982 13920 30006 14160
rect 30242 13920 30246 14160
rect 30266 13920 30302 14160
rect 33982 14160 34302 14222
rect 29982 13896 30302 13920
rect 32366 13916 32606 13940
rect 32366 13740 32390 13916
rect 32582 13740 32606 13916
rect 33982 13920 34006 14160
rect 34242 13920 34246 14160
rect 34266 13920 34302 14160
rect 37982 14160 38302 14222
rect 33982 13896 34302 13920
rect 36366 13916 36606 13940
rect 36366 13740 36390 13916
rect 36582 13740 36606 13916
rect 37982 13920 38006 14160
rect 38242 13920 38246 14160
rect 38266 13920 38302 14160
rect 37982 13896 38302 13920
use fgcell_amp_MOS_cap_thick_poly  fgcell_amp_MOS_cap_thick_poly_0
array 0 9 4000 0 4 3000
timestamp 1717597427
transform 1 0 -140 0 1 22210
box 74 -7210 4106 -4964
use fgcell_amp_MOS_cap_thin_poly  fgcell_amp_MOS_cap_thin_poly_0
array 0 9 4000 0 4 3000
timestamp 1717597427
transform 1 0 -140 0 1 7210
box 74 -7210 4106 -4964
<< end >>
