magic
tech sky130A
timestamp 1716502360
<< nwell >>
rect 10 860 570 1450
<< mvnmos >>
rect 100 600 200 750
rect 250 600 350 750
rect 100 350 200 500
rect 250 350 350 500
rect 100 100 200 250
rect 250 100 350 250
<< mvpmos >>
rect 100 1200 200 1350
rect 250 1200 350 1350
rect 100 900 200 1050
rect 250 900 350 1050
<< mvndiff >>
rect 50 740 100 750
rect 50 610 60 740
rect 90 610 100 740
rect 50 600 100 610
rect 200 740 250 750
rect 200 610 210 740
rect 240 610 250 740
rect 200 600 250 610
rect 350 740 400 750
rect 350 610 360 740
rect 390 610 400 740
rect 350 600 400 610
rect 50 490 100 500
rect 50 360 60 490
rect 90 360 100 490
rect 50 350 100 360
rect 200 350 250 500
rect 350 490 400 500
rect 350 360 360 490
rect 390 360 400 490
rect 350 350 400 360
rect 50 240 100 250
rect 50 110 60 240
rect 90 110 100 240
rect 50 100 100 110
rect 200 240 250 250
rect 200 110 210 240
rect 240 110 250 240
rect 200 100 250 110
rect 350 240 400 250
rect 350 110 360 240
rect 390 110 400 240
rect 350 100 400 110
<< mvpdiff >>
rect 50 1340 100 1350
rect 50 1210 60 1340
rect 90 1210 100 1340
rect 50 1200 100 1210
rect 200 1340 250 1350
rect 200 1210 210 1340
rect 240 1210 250 1340
rect 200 1200 250 1210
rect 350 1340 400 1350
rect 350 1210 360 1340
rect 390 1210 400 1340
rect 350 1200 400 1210
rect 50 1040 100 1050
rect 50 910 60 1040
rect 90 910 100 1040
rect 50 900 100 910
rect 200 1040 250 1050
rect 200 910 210 1040
rect 240 910 250 1040
rect 200 900 250 910
rect 350 1040 400 1050
rect 350 910 360 1040
rect 390 910 400 1040
rect 350 900 400 910
<< mvndiffc >>
rect 60 610 90 740
rect 210 610 240 740
rect 360 610 390 740
rect 60 360 90 490
rect 360 360 390 490
rect 60 110 90 240
rect 210 110 240 240
rect 360 110 390 240
<< mvpdiffc >>
rect 60 1210 90 1340
rect 210 1210 240 1340
rect 360 1210 390 1340
rect 60 910 90 1040
rect 210 910 240 1040
rect 360 910 390 1040
<< mvpsubdiff >>
rect 470 480 530 500
rect 470 370 490 480
rect 510 370 530 480
rect 470 350 530 370
<< mvnsubdiff >>
rect 470 1340 530 1350
rect 470 1210 490 1340
rect 510 1210 530 1340
rect 470 1200 530 1210
<< mvpsubdiffcont >>
rect 490 370 510 480
<< mvnsubdiffcont >>
rect 490 1210 510 1340
<< poly >>
rect 100 1350 200 1370
rect 250 1350 350 1370
rect 100 1180 200 1200
rect 250 1180 350 1200
rect 100 1170 350 1180
rect 100 1150 260 1170
rect 340 1150 350 1170
rect 100 1140 350 1150
rect 100 1050 200 1070
rect 250 1050 350 1070
rect 100 880 200 900
rect 250 880 350 900
rect 100 870 350 880
rect 100 850 110 870
rect 190 850 350 870
rect 100 840 350 850
rect 100 790 200 800
rect 100 770 110 790
rect 190 770 200 790
rect 100 750 200 770
rect 250 790 350 800
rect 250 770 260 790
rect 340 770 350 790
rect 250 750 350 770
rect 100 580 200 600
rect 250 580 350 600
rect 100 500 200 520
rect 250 500 350 520
rect 100 340 200 350
rect 250 340 350 350
rect 100 330 350 340
rect 100 310 110 330
rect 190 310 350 330
rect 100 300 350 310
rect 100 250 200 270
rect 250 250 350 270
rect 100 90 200 100
rect 250 90 350 100
rect 100 80 350 90
rect 100 40 110 80
rect 190 40 350 80
rect 100 30 350 40
<< polycont >>
rect 260 1150 340 1170
rect 110 850 190 870
rect 110 770 190 790
rect 260 770 340 790
rect 110 310 190 330
rect 110 40 190 80
<< locali >>
rect 60 1340 90 1350
rect 0 1240 60 1250
rect 0 1210 10 1240
rect 40 1210 60 1240
rect 0 1200 90 1210
rect 210 1340 240 1350
rect 60 1040 90 1050
rect 60 880 90 910
rect 210 1040 240 1210
rect 360 1340 410 1350
rect 390 1210 410 1340
rect 360 1180 410 1210
rect 490 1340 510 1350
rect 490 1200 510 1210
rect 260 1170 410 1180
rect 340 1150 370 1170
rect 260 1140 370 1150
rect 400 1140 410 1170
rect 260 1130 410 1140
rect 210 900 240 910
rect 360 1040 530 1050
rect 390 910 490 1040
rect 520 910 530 1040
rect 360 900 530 910
rect 60 870 200 880
rect 60 850 110 870
rect 190 850 200 870
rect 60 840 200 850
rect 60 740 90 840
rect 110 790 190 800
rect 110 760 190 770
rect 260 790 340 800
rect 260 760 340 770
rect 60 600 90 610
rect 210 740 240 750
rect 210 570 240 610
rect 360 740 450 750
rect 390 710 410 740
rect 440 710 450 740
rect 390 700 450 710
rect 360 600 390 610
rect 60 530 240 570
rect 60 490 90 530
rect 60 350 90 360
rect 360 490 530 500
rect 390 480 530 490
rect 390 370 490 480
rect 510 370 530 480
rect 390 360 530 370
rect 360 350 530 360
rect 110 330 190 340
rect 110 300 190 310
rect 0 240 90 250
rect 0 210 10 240
rect 40 210 60 240
rect 0 200 60 210
rect 60 80 90 110
rect 210 240 240 250
rect 210 100 240 110
rect 360 240 450 250
rect 390 210 410 240
rect 440 210 450 240
rect 390 200 450 210
rect 360 100 390 110
rect 60 40 110 80
rect 190 40 200 80
<< viali >>
rect 10 1210 40 1240
rect 370 1140 400 1170
rect 210 910 240 1040
rect 490 910 520 1040
rect 410 710 440 740
rect 10 210 40 240
rect 210 110 240 240
rect 410 210 440 240
<< metal1 >>
rect 0 1240 50 1250
rect 0 1210 10 1240
rect 40 1210 50 1240
rect 0 240 50 1210
rect 200 1040 250 1350
rect 360 1170 450 1180
rect 360 1140 370 1170
rect 400 1140 450 1170
rect 360 1130 450 1140
rect 200 910 210 1040
rect 240 910 250 1040
rect 200 900 250 910
rect 400 740 450 1130
rect 400 710 410 740
rect 440 710 450 740
rect 400 700 450 710
rect 480 1040 530 1050
rect 480 910 490 1040
rect 520 910 530 1040
rect 480 580 530 910
rect 400 530 530 580
rect 0 210 10 240
rect 40 210 50 240
rect 0 200 50 210
rect 200 240 250 250
rect 200 110 210 240
rect 240 150 250 240
rect 400 240 450 530
rect 400 210 410 240
rect 440 210 450 240
rect 400 200 450 210
rect 240 110 530 150
rect 200 100 530 110
<< end >>
