magic
tech sky130A
magscale 1 2
timestamp 1717582298
<< dnwell >>
rect 618 14749 14328 36195
<< nwell >>
rect 509 35931 14439 36306
rect 509 15013 824 35931
rect 1585 28325 13415 28988
rect 1585 27635 2328 28325
rect 12672 27635 13415 28325
rect 1585 26891 13415 27635
rect 2320 25375 12656 26045
rect 14064 15013 14439 35931
rect 509 14638 14439 15013
<< pwell >>
rect 211 36376 14742 36613
rect 211 14567 448 36376
rect 1085 34590 13905 34760
rect 1085 15358 1255 34590
rect 2338 27645 12662 28315
rect 1722 26165 13254 26611
rect 1722 25255 2168 26165
rect 12808 25255 13254 26165
rect 1722 24809 13254 25255
rect 13735 15358 13905 34590
rect 1085 15188 13905 15358
rect 14505 14567 14742 36376
rect 211 14330 14742 14567
<< mvpsubdiff >>
rect 237 36510 14716 36587
rect 237 36476 447 36510
rect 481 36476 515 36510
rect 549 36476 583 36510
rect 617 36476 651 36510
rect 685 36476 719 36510
rect 753 36476 787 36510
rect 821 36476 855 36510
rect 889 36476 923 36510
rect 957 36476 991 36510
rect 1025 36476 1059 36510
rect 1093 36476 1127 36510
rect 1161 36476 1195 36510
rect 1229 36476 1263 36510
rect 1297 36476 1331 36510
rect 1365 36476 1399 36510
rect 1433 36476 1467 36510
rect 1501 36476 1535 36510
rect 1569 36476 1603 36510
rect 1637 36476 1671 36510
rect 1705 36476 1739 36510
rect 1773 36476 1807 36510
rect 1841 36476 1875 36510
rect 1909 36476 1943 36510
rect 1977 36476 2011 36510
rect 2045 36476 2079 36510
rect 2113 36476 2147 36510
rect 2181 36476 2215 36510
rect 2249 36476 2283 36510
rect 2317 36476 2351 36510
rect 2385 36476 2419 36510
rect 2453 36476 2487 36510
rect 2521 36476 2555 36510
rect 2589 36476 2623 36510
rect 2657 36476 2691 36510
rect 2725 36476 2759 36510
rect 2793 36476 2827 36510
rect 2861 36476 2895 36510
rect 2929 36476 2963 36510
rect 2997 36476 3031 36510
rect 3065 36476 3099 36510
rect 3133 36476 3167 36510
rect 3201 36476 3235 36510
rect 3269 36476 3303 36510
rect 3337 36476 3371 36510
rect 3405 36476 3439 36510
rect 3473 36476 3507 36510
rect 3541 36476 3575 36510
rect 3609 36476 3643 36510
rect 3677 36476 3711 36510
rect 3745 36476 3779 36510
rect 3813 36476 3847 36510
rect 3881 36476 3915 36510
rect 3949 36476 3983 36510
rect 4017 36476 4051 36510
rect 4085 36476 4119 36510
rect 4153 36476 4187 36510
rect 4221 36476 4255 36510
rect 4289 36476 4323 36510
rect 4357 36476 4391 36510
rect 4425 36476 4459 36510
rect 4493 36476 4527 36510
rect 4561 36476 4595 36510
rect 4629 36476 4663 36510
rect 4697 36476 4731 36510
rect 4765 36476 4799 36510
rect 4833 36476 4867 36510
rect 4901 36476 4935 36510
rect 4969 36476 5003 36510
rect 5037 36476 5071 36510
rect 5105 36476 5139 36510
rect 5173 36476 5207 36510
rect 5241 36476 5275 36510
rect 5309 36476 5343 36510
rect 5377 36476 5411 36510
rect 5445 36476 5479 36510
rect 5513 36476 5547 36510
rect 5581 36476 5615 36510
rect 5649 36476 5683 36510
rect 5717 36476 5751 36510
rect 5785 36476 5819 36510
rect 5853 36476 5887 36510
rect 5921 36476 5955 36510
rect 5989 36476 6023 36510
rect 6057 36476 6091 36510
rect 6125 36476 6159 36510
rect 6193 36476 6227 36510
rect 6261 36476 6295 36510
rect 6329 36476 6363 36510
rect 6397 36476 6431 36510
rect 6465 36476 6499 36510
rect 6533 36476 6567 36510
rect 6601 36476 6635 36510
rect 6669 36476 6703 36510
rect 6737 36476 6771 36510
rect 6805 36476 6839 36510
rect 6873 36476 6907 36510
rect 6941 36476 6975 36510
rect 7009 36476 7043 36510
rect 7077 36476 7111 36510
rect 7145 36476 7179 36510
rect 7213 36476 7247 36510
rect 7281 36476 7315 36510
rect 7349 36476 7383 36510
rect 7417 36476 7451 36510
rect 7485 36476 7519 36510
rect 7553 36476 7587 36510
rect 7621 36476 7655 36510
rect 7689 36476 7723 36510
rect 7757 36476 7791 36510
rect 7825 36476 7859 36510
rect 7893 36476 7927 36510
rect 7961 36476 7995 36510
rect 8029 36476 8063 36510
rect 8097 36476 8131 36510
rect 8165 36476 8199 36510
rect 8233 36476 8267 36510
rect 8301 36476 8335 36510
rect 8369 36476 8403 36510
rect 8437 36476 8471 36510
rect 8505 36476 8539 36510
rect 8573 36476 8607 36510
rect 8641 36476 8675 36510
rect 8709 36476 8743 36510
rect 8777 36476 8811 36510
rect 8845 36476 8879 36510
rect 8913 36476 8947 36510
rect 8981 36476 9015 36510
rect 9049 36476 9083 36510
rect 9117 36476 9151 36510
rect 9185 36476 9219 36510
rect 9253 36476 9287 36510
rect 9321 36476 9355 36510
rect 9389 36476 9423 36510
rect 9457 36476 9491 36510
rect 9525 36476 9559 36510
rect 9593 36476 9627 36510
rect 9661 36476 9695 36510
rect 9729 36476 9763 36510
rect 9797 36476 9831 36510
rect 9865 36476 9899 36510
rect 9933 36476 9967 36510
rect 10001 36476 10035 36510
rect 10069 36476 10103 36510
rect 10137 36476 10171 36510
rect 10205 36476 10239 36510
rect 10273 36476 10307 36510
rect 10341 36476 10375 36510
rect 10409 36476 10443 36510
rect 10477 36476 10511 36510
rect 10545 36476 10579 36510
rect 10613 36476 10647 36510
rect 10681 36476 10715 36510
rect 10749 36476 10783 36510
rect 10817 36476 10851 36510
rect 10885 36476 10919 36510
rect 10953 36476 10987 36510
rect 11021 36476 11055 36510
rect 11089 36476 11123 36510
rect 11157 36476 11191 36510
rect 11225 36476 11259 36510
rect 11293 36476 11327 36510
rect 11361 36476 11395 36510
rect 11429 36476 11463 36510
rect 11497 36476 11531 36510
rect 11565 36476 11599 36510
rect 11633 36476 11667 36510
rect 11701 36476 11735 36510
rect 11769 36476 11803 36510
rect 11837 36476 11871 36510
rect 11905 36476 11939 36510
rect 11973 36476 12007 36510
rect 12041 36476 12075 36510
rect 12109 36476 12143 36510
rect 12177 36476 12211 36510
rect 12245 36476 12279 36510
rect 12313 36476 12347 36510
rect 12381 36476 12415 36510
rect 12449 36476 12483 36510
rect 12517 36476 12551 36510
rect 12585 36476 12619 36510
rect 12653 36476 12687 36510
rect 12721 36476 12755 36510
rect 12789 36476 12823 36510
rect 12857 36476 12891 36510
rect 12925 36476 12959 36510
rect 12993 36476 13027 36510
rect 13061 36476 13095 36510
rect 13129 36476 13163 36510
rect 13197 36476 13231 36510
rect 13265 36476 13299 36510
rect 13333 36476 13367 36510
rect 13401 36476 13435 36510
rect 13469 36476 13503 36510
rect 13537 36476 13571 36510
rect 13605 36476 13639 36510
rect 13673 36476 13707 36510
rect 13741 36476 13775 36510
rect 13809 36476 13843 36510
rect 13877 36476 13911 36510
rect 13945 36476 13979 36510
rect 14013 36476 14047 36510
rect 14081 36476 14115 36510
rect 14149 36476 14183 36510
rect 14217 36476 14251 36510
rect 14285 36476 14319 36510
rect 14353 36476 14387 36510
rect 14421 36476 14455 36510
rect 14489 36476 14716 36510
rect 237 36402 14716 36476
rect 237 36369 422 36402
rect 237 36335 304 36369
rect 338 36335 422 36369
rect 237 36301 422 36335
rect 237 36267 304 36301
rect 338 36267 422 36301
rect 237 36233 422 36267
rect 14531 36375 14716 36402
rect 14531 36341 14599 36375
rect 14633 36341 14716 36375
rect 14531 36307 14716 36341
rect 14531 36273 14599 36307
rect 14633 36273 14716 36307
rect 237 36199 304 36233
rect 338 36199 422 36233
rect 237 36165 422 36199
rect 237 36131 304 36165
rect 338 36131 422 36165
rect 237 36097 422 36131
rect 237 36063 304 36097
rect 338 36063 422 36097
rect 237 36029 422 36063
rect 237 35995 304 36029
rect 338 35995 422 36029
rect 237 35961 422 35995
rect 237 35927 304 35961
rect 338 35927 422 35961
rect 237 35893 422 35927
rect 237 35859 304 35893
rect 338 35859 422 35893
rect 237 35825 422 35859
rect 237 35791 304 35825
rect 338 35791 422 35825
rect 237 35757 422 35791
rect 237 35723 304 35757
rect 338 35723 422 35757
rect 237 35689 422 35723
rect 237 35655 304 35689
rect 338 35655 422 35689
rect 237 35621 422 35655
rect 237 35587 304 35621
rect 338 35587 422 35621
rect 237 35553 422 35587
rect 237 35519 304 35553
rect 338 35519 422 35553
rect 237 35485 422 35519
rect 237 35451 304 35485
rect 338 35451 422 35485
rect 237 35417 422 35451
rect 237 35383 304 35417
rect 338 35383 422 35417
rect 237 35349 422 35383
rect 237 35315 304 35349
rect 338 35315 422 35349
rect 237 35281 422 35315
rect 237 35247 304 35281
rect 338 35247 422 35281
rect 237 35213 422 35247
rect 237 35179 304 35213
rect 338 35179 422 35213
rect 237 35145 422 35179
rect 237 35111 304 35145
rect 338 35111 422 35145
rect 237 35077 422 35111
rect 237 35043 304 35077
rect 338 35043 422 35077
rect 237 35009 422 35043
rect 237 34975 304 35009
rect 338 34975 422 35009
rect 237 34941 422 34975
rect 237 34907 304 34941
rect 338 34907 422 34941
rect 237 34873 422 34907
rect 237 34839 304 34873
rect 338 34839 422 34873
rect 237 34805 422 34839
rect 237 34771 304 34805
rect 338 34771 422 34805
rect 237 34737 422 34771
rect 237 34703 304 34737
rect 338 34703 422 34737
rect 237 34669 422 34703
rect 237 34635 304 34669
rect 338 34635 422 34669
rect 237 34601 422 34635
rect 237 34567 304 34601
rect 338 34567 422 34601
rect 237 34533 422 34567
rect 237 34499 304 34533
rect 338 34499 422 34533
rect 237 34465 422 34499
rect 237 34431 304 34465
rect 338 34431 422 34465
rect 237 34397 422 34431
rect 237 34363 304 34397
rect 338 34363 422 34397
rect 237 34329 422 34363
rect 237 34295 304 34329
rect 338 34295 422 34329
rect 237 34261 422 34295
rect 237 34227 304 34261
rect 338 34227 422 34261
rect 237 34193 422 34227
rect 237 34159 304 34193
rect 338 34159 422 34193
rect 237 34125 422 34159
rect 237 34091 304 34125
rect 338 34091 422 34125
rect 237 34057 422 34091
rect 237 34023 304 34057
rect 338 34023 422 34057
rect 237 33989 422 34023
rect 237 33955 304 33989
rect 338 33955 422 33989
rect 237 33921 422 33955
rect 237 33887 304 33921
rect 338 33887 422 33921
rect 237 33853 422 33887
rect 237 33819 304 33853
rect 338 33819 422 33853
rect 237 33785 422 33819
rect 237 33751 304 33785
rect 338 33751 422 33785
rect 237 33717 422 33751
rect 237 33683 304 33717
rect 338 33683 422 33717
rect 237 33649 422 33683
rect 237 33615 304 33649
rect 338 33615 422 33649
rect 237 33581 422 33615
rect 237 33547 304 33581
rect 338 33547 422 33581
rect 237 33513 422 33547
rect 237 33479 304 33513
rect 338 33479 422 33513
rect 237 33445 422 33479
rect 237 33411 304 33445
rect 338 33411 422 33445
rect 237 33377 422 33411
rect 237 33343 304 33377
rect 338 33343 422 33377
rect 237 33309 422 33343
rect 237 33275 304 33309
rect 338 33275 422 33309
rect 237 33241 422 33275
rect 237 33207 304 33241
rect 338 33207 422 33241
rect 237 33173 422 33207
rect 237 33139 304 33173
rect 338 33139 422 33173
rect 237 33105 422 33139
rect 237 33071 304 33105
rect 338 33071 422 33105
rect 237 33037 422 33071
rect 237 33003 304 33037
rect 338 33003 422 33037
rect 237 32969 422 33003
rect 237 32935 304 32969
rect 338 32935 422 32969
rect 237 32901 422 32935
rect 237 32867 304 32901
rect 338 32867 422 32901
rect 237 32833 422 32867
rect 237 32799 304 32833
rect 338 32799 422 32833
rect 237 32765 422 32799
rect 237 32731 304 32765
rect 338 32731 422 32765
rect 237 32697 422 32731
rect 237 32663 304 32697
rect 338 32663 422 32697
rect 237 32629 422 32663
rect 237 32595 304 32629
rect 338 32595 422 32629
rect 237 32561 422 32595
rect 237 32527 304 32561
rect 338 32527 422 32561
rect 237 32493 422 32527
rect 237 32459 304 32493
rect 338 32459 422 32493
rect 237 32425 422 32459
rect 237 32391 304 32425
rect 338 32391 422 32425
rect 237 32357 422 32391
rect 237 32323 304 32357
rect 338 32323 422 32357
rect 237 32289 422 32323
rect 237 32255 304 32289
rect 338 32255 422 32289
rect 237 32221 422 32255
rect 237 32187 304 32221
rect 338 32187 422 32221
rect 237 32153 422 32187
rect 237 32119 304 32153
rect 338 32119 422 32153
rect 237 32085 422 32119
rect 237 32051 304 32085
rect 338 32051 422 32085
rect 237 32017 422 32051
rect 237 31983 304 32017
rect 338 31983 422 32017
rect 237 31949 422 31983
rect 237 31915 304 31949
rect 338 31915 422 31949
rect 237 31881 422 31915
rect 237 31847 304 31881
rect 338 31847 422 31881
rect 237 31813 422 31847
rect 237 31779 304 31813
rect 338 31779 422 31813
rect 237 31745 422 31779
rect 237 31711 304 31745
rect 338 31711 422 31745
rect 237 31677 422 31711
rect 237 31643 304 31677
rect 338 31643 422 31677
rect 237 31609 422 31643
rect 237 31575 304 31609
rect 338 31575 422 31609
rect 237 31541 422 31575
rect 237 31507 304 31541
rect 338 31507 422 31541
rect 237 31473 422 31507
rect 237 31439 304 31473
rect 338 31439 422 31473
rect 237 31405 422 31439
rect 237 31371 304 31405
rect 338 31371 422 31405
rect 237 31337 422 31371
rect 237 31303 304 31337
rect 338 31303 422 31337
rect 237 31269 422 31303
rect 237 31235 304 31269
rect 338 31235 422 31269
rect 237 31201 422 31235
rect 237 31167 304 31201
rect 338 31167 422 31201
rect 237 31133 422 31167
rect 237 31099 304 31133
rect 338 31099 422 31133
rect 237 31065 422 31099
rect 237 31031 304 31065
rect 338 31031 422 31065
rect 237 30997 422 31031
rect 237 30963 304 30997
rect 338 30963 422 30997
rect 237 30929 422 30963
rect 237 30895 304 30929
rect 338 30895 422 30929
rect 237 30861 422 30895
rect 237 30827 304 30861
rect 338 30827 422 30861
rect 237 30793 422 30827
rect 237 30759 304 30793
rect 338 30759 422 30793
rect 237 30725 422 30759
rect 237 30691 304 30725
rect 338 30691 422 30725
rect 237 30657 422 30691
rect 237 30623 304 30657
rect 338 30623 422 30657
rect 237 30589 422 30623
rect 237 30555 304 30589
rect 338 30555 422 30589
rect 237 30521 422 30555
rect 237 30487 304 30521
rect 338 30487 422 30521
rect 237 30453 422 30487
rect 237 30419 304 30453
rect 338 30419 422 30453
rect 237 30385 422 30419
rect 237 30351 304 30385
rect 338 30351 422 30385
rect 237 30317 422 30351
rect 237 30283 304 30317
rect 338 30283 422 30317
rect 237 30249 422 30283
rect 237 30215 304 30249
rect 338 30215 422 30249
rect 237 30181 422 30215
rect 237 30147 304 30181
rect 338 30147 422 30181
rect 237 30113 422 30147
rect 237 30079 304 30113
rect 338 30079 422 30113
rect 237 30045 422 30079
rect 237 30011 304 30045
rect 338 30011 422 30045
rect 237 29977 422 30011
rect 237 29943 304 29977
rect 338 29943 422 29977
rect 237 29909 422 29943
rect 237 29875 304 29909
rect 338 29875 422 29909
rect 237 29841 422 29875
rect 237 29807 304 29841
rect 338 29807 422 29841
rect 237 29773 422 29807
rect 237 29739 304 29773
rect 338 29739 422 29773
rect 237 29705 422 29739
rect 237 29671 304 29705
rect 338 29671 422 29705
rect 237 29637 422 29671
rect 237 29603 304 29637
rect 338 29603 422 29637
rect 237 29569 422 29603
rect 237 29535 304 29569
rect 338 29535 422 29569
rect 237 29501 422 29535
rect 237 29467 304 29501
rect 338 29467 422 29501
rect 237 29433 422 29467
rect 237 29399 304 29433
rect 338 29399 422 29433
rect 237 29365 422 29399
rect 237 29331 304 29365
rect 338 29331 422 29365
rect 237 29297 422 29331
rect 237 29263 304 29297
rect 338 29263 422 29297
rect 237 29229 422 29263
rect 237 29195 304 29229
rect 338 29195 422 29229
rect 237 29161 422 29195
rect 237 29127 304 29161
rect 338 29127 422 29161
rect 237 29093 422 29127
rect 237 29059 304 29093
rect 338 29059 422 29093
rect 237 29025 422 29059
rect 237 28991 304 29025
rect 338 28991 422 29025
rect 237 28957 422 28991
rect 237 28923 304 28957
rect 338 28923 422 28957
rect 237 28889 422 28923
rect 237 28855 304 28889
rect 338 28855 422 28889
rect 237 28821 422 28855
rect 237 28787 304 28821
rect 338 28787 422 28821
rect 237 28753 422 28787
rect 237 28719 304 28753
rect 338 28719 422 28753
rect 237 28685 422 28719
rect 237 28651 304 28685
rect 338 28651 422 28685
rect 237 28617 422 28651
rect 237 28583 304 28617
rect 338 28583 422 28617
rect 237 28549 422 28583
rect 237 28515 304 28549
rect 338 28515 422 28549
rect 237 28481 422 28515
rect 237 28447 304 28481
rect 338 28447 422 28481
rect 237 28413 422 28447
rect 237 28379 304 28413
rect 338 28379 422 28413
rect 237 28345 422 28379
rect 237 28311 304 28345
rect 338 28311 422 28345
rect 237 28277 422 28311
rect 237 28243 304 28277
rect 338 28243 422 28277
rect 237 28209 422 28243
rect 237 28175 304 28209
rect 338 28175 422 28209
rect 237 28141 422 28175
rect 237 28107 304 28141
rect 338 28107 422 28141
rect 237 28073 422 28107
rect 237 28039 304 28073
rect 338 28039 422 28073
rect 237 28005 422 28039
rect 237 27971 304 28005
rect 338 27971 422 28005
rect 237 27937 422 27971
rect 237 27903 304 27937
rect 338 27903 422 27937
rect 237 27869 422 27903
rect 237 27835 304 27869
rect 338 27835 422 27869
rect 237 27801 422 27835
rect 237 27767 304 27801
rect 338 27767 422 27801
rect 237 27733 422 27767
rect 237 27699 304 27733
rect 338 27699 422 27733
rect 237 27665 422 27699
rect 237 27631 304 27665
rect 338 27631 422 27665
rect 237 27597 422 27631
rect 237 27563 304 27597
rect 338 27563 422 27597
rect 237 27529 422 27563
rect 237 27495 304 27529
rect 338 27495 422 27529
rect 237 27461 422 27495
rect 237 27427 304 27461
rect 338 27427 422 27461
rect 237 27393 422 27427
rect 237 27359 304 27393
rect 338 27359 422 27393
rect 237 27325 422 27359
rect 237 27291 304 27325
rect 338 27291 422 27325
rect 237 27257 422 27291
rect 237 27223 304 27257
rect 338 27223 422 27257
rect 237 27189 422 27223
rect 237 27155 304 27189
rect 338 27155 422 27189
rect 237 27121 422 27155
rect 237 27087 304 27121
rect 338 27087 422 27121
rect 237 27053 422 27087
rect 237 27019 304 27053
rect 338 27019 422 27053
rect 237 26985 422 27019
rect 237 26951 304 26985
rect 338 26951 422 26985
rect 237 26917 422 26951
rect 237 26883 304 26917
rect 338 26883 422 26917
rect 237 26849 422 26883
rect 237 26815 304 26849
rect 338 26815 422 26849
rect 237 26781 422 26815
rect 237 26747 304 26781
rect 338 26747 422 26781
rect 237 26713 422 26747
rect 237 26679 304 26713
rect 338 26679 422 26713
rect 237 26645 422 26679
rect 237 26611 304 26645
rect 338 26611 422 26645
rect 237 26577 422 26611
rect 237 26543 304 26577
rect 338 26543 422 26577
rect 237 26509 422 26543
rect 237 26475 304 26509
rect 338 26475 422 26509
rect 237 26441 422 26475
rect 237 26407 304 26441
rect 338 26407 422 26441
rect 237 26373 422 26407
rect 237 26339 304 26373
rect 338 26339 422 26373
rect 237 26305 422 26339
rect 237 26271 304 26305
rect 338 26271 422 26305
rect 237 26237 422 26271
rect 237 26203 304 26237
rect 338 26203 422 26237
rect 237 26169 422 26203
rect 237 26135 304 26169
rect 338 26135 422 26169
rect 237 26101 422 26135
rect 237 26067 304 26101
rect 338 26067 422 26101
rect 237 26033 422 26067
rect 237 25999 304 26033
rect 338 25999 422 26033
rect 237 25965 422 25999
rect 237 25931 304 25965
rect 338 25931 422 25965
rect 237 25897 422 25931
rect 237 25863 304 25897
rect 338 25863 422 25897
rect 237 25829 422 25863
rect 237 25795 304 25829
rect 338 25795 422 25829
rect 237 25761 422 25795
rect 237 25727 304 25761
rect 338 25727 422 25761
rect 237 25693 422 25727
rect 237 25659 304 25693
rect 338 25659 422 25693
rect 237 25625 422 25659
rect 237 25591 304 25625
rect 338 25591 422 25625
rect 237 25557 422 25591
rect 237 25523 304 25557
rect 338 25523 422 25557
rect 237 25489 422 25523
rect 237 25455 304 25489
rect 338 25455 422 25489
rect 237 25421 422 25455
rect 237 25387 304 25421
rect 338 25387 422 25421
rect 237 25353 422 25387
rect 237 25319 304 25353
rect 338 25319 422 25353
rect 237 25285 422 25319
rect 237 25251 304 25285
rect 338 25251 422 25285
rect 237 25217 422 25251
rect 237 25183 304 25217
rect 338 25183 422 25217
rect 237 25149 422 25183
rect 237 25115 304 25149
rect 338 25115 422 25149
rect 237 25081 422 25115
rect 237 25047 304 25081
rect 338 25047 422 25081
rect 237 25013 422 25047
rect 237 24979 304 25013
rect 338 24979 422 25013
rect 237 24945 422 24979
rect 237 24911 304 24945
rect 338 24911 422 24945
rect 237 24877 422 24911
rect 237 24843 304 24877
rect 338 24843 422 24877
rect 237 24809 422 24843
rect 237 24775 304 24809
rect 338 24775 422 24809
rect 237 24741 422 24775
rect 237 24707 304 24741
rect 338 24707 422 24741
rect 237 24673 422 24707
rect 237 24639 304 24673
rect 338 24639 422 24673
rect 237 24605 422 24639
rect 237 24571 304 24605
rect 338 24571 422 24605
rect 237 24537 422 24571
rect 237 24503 304 24537
rect 338 24503 422 24537
rect 237 24469 422 24503
rect 237 24435 304 24469
rect 338 24435 422 24469
rect 237 24401 422 24435
rect 237 24367 304 24401
rect 338 24367 422 24401
rect 237 24333 422 24367
rect 237 24299 304 24333
rect 338 24299 422 24333
rect 237 24265 422 24299
rect 237 24231 304 24265
rect 338 24231 422 24265
rect 237 24197 422 24231
rect 237 24163 304 24197
rect 338 24163 422 24197
rect 237 24129 422 24163
rect 237 24095 304 24129
rect 338 24095 422 24129
rect 237 24061 422 24095
rect 237 24027 304 24061
rect 338 24027 422 24061
rect 237 23993 422 24027
rect 237 23959 304 23993
rect 338 23959 422 23993
rect 237 23925 422 23959
rect 237 23891 304 23925
rect 338 23891 422 23925
rect 237 23857 422 23891
rect 237 23823 304 23857
rect 338 23823 422 23857
rect 237 23789 422 23823
rect 237 23755 304 23789
rect 338 23755 422 23789
rect 237 23721 422 23755
rect 237 23687 304 23721
rect 338 23687 422 23721
rect 237 23653 422 23687
rect 237 23619 304 23653
rect 338 23619 422 23653
rect 237 23585 422 23619
rect 237 23551 304 23585
rect 338 23551 422 23585
rect 237 23517 422 23551
rect 237 23483 304 23517
rect 338 23483 422 23517
rect 237 23449 422 23483
rect 237 23415 304 23449
rect 338 23415 422 23449
rect 237 23381 422 23415
rect 237 23347 304 23381
rect 338 23347 422 23381
rect 237 23313 422 23347
rect 237 23279 304 23313
rect 338 23279 422 23313
rect 237 23245 422 23279
rect 237 23211 304 23245
rect 338 23211 422 23245
rect 237 23177 422 23211
rect 237 23143 304 23177
rect 338 23143 422 23177
rect 237 23109 422 23143
rect 237 23075 304 23109
rect 338 23075 422 23109
rect 237 23041 422 23075
rect 237 23007 304 23041
rect 338 23007 422 23041
rect 237 22973 422 23007
rect 237 22939 304 22973
rect 338 22939 422 22973
rect 237 22905 422 22939
rect 237 22871 304 22905
rect 338 22871 422 22905
rect 237 22837 422 22871
rect 237 22803 304 22837
rect 338 22803 422 22837
rect 237 22769 422 22803
rect 237 22735 304 22769
rect 338 22735 422 22769
rect 237 22701 422 22735
rect 237 22667 304 22701
rect 338 22667 422 22701
rect 237 22633 422 22667
rect 237 22599 304 22633
rect 338 22599 422 22633
rect 237 22565 422 22599
rect 237 22531 304 22565
rect 338 22531 422 22565
rect 237 22497 422 22531
rect 237 22463 304 22497
rect 338 22463 422 22497
rect 237 22429 422 22463
rect 237 22395 304 22429
rect 338 22395 422 22429
rect 237 22361 422 22395
rect 237 22327 304 22361
rect 338 22327 422 22361
rect 237 22293 422 22327
rect 237 22259 304 22293
rect 338 22259 422 22293
rect 237 22225 422 22259
rect 237 22191 304 22225
rect 338 22191 422 22225
rect 237 22157 422 22191
rect 237 22123 304 22157
rect 338 22123 422 22157
rect 237 22089 422 22123
rect 237 22055 304 22089
rect 338 22055 422 22089
rect 237 22021 422 22055
rect 237 21987 304 22021
rect 338 21987 422 22021
rect 237 21953 422 21987
rect 237 21919 304 21953
rect 338 21919 422 21953
rect 237 21885 422 21919
rect 237 21851 304 21885
rect 338 21851 422 21885
rect 237 21817 422 21851
rect 237 21783 304 21817
rect 338 21783 422 21817
rect 237 21749 422 21783
rect 237 21715 304 21749
rect 338 21715 422 21749
rect 237 21681 422 21715
rect 237 21647 304 21681
rect 338 21647 422 21681
rect 237 21613 422 21647
rect 237 21579 304 21613
rect 338 21579 422 21613
rect 237 21545 422 21579
rect 237 21511 304 21545
rect 338 21511 422 21545
rect 237 21477 422 21511
rect 237 21443 304 21477
rect 338 21443 422 21477
rect 237 21409 422 21443
rect 237 21375 304 21409
rect 338 21375 422 21409
rect 237 21341 422 21375
rect 237 21307 304 21341
rect 338 21307 422 21341
rect 237 21273 422 21307
rect 237 21239 304 21273
rect 338 21239 422 21273
rect 237 21205 422 21239
rect 237 21171 304 21205
rect 338 21171 422 21205
rect 237 21137 422 21171
rect 237 21103 304 21137
rect 338 21103 422 21137
rect 237 21069 422 21103
rect 237 21035 304 21069
rect 338 21035 422 21069
rect 237 21001 422 21035
rect 237 20967 304 21001
rect 338 20967 422 21001
rect 237 20933 422 20967
rect 237 20899 304 20933
rect 338 20899 422 20933
rect 237 20865 422 20899
rect 237 20831 304 20865
rect 338 20831 422 20865
rect 237 20797 422 20831
rect 237 20763 304 20797
rect 338 20763 422 20797
rect 237 20729 422 20763
rect 237 20695 304 20729
rect 338 20695 422 20729
rect 237 20661 422 20695
rect 237 20627 304 20661
rect 338 20627 422 20661
rect 237 20593 422 20627
rect 237 20559 304 20593
rect 338 20559 422 20593
rect 237 20525 422 20559
rect 237 20491 304 20525
rect 338 20491 422 20525
rect 237 20457 422 20491
rect 237 20423 304 20457
rect 338 20423 422 20457
rect 237 20389 422 20423
rect 237 20355 304 20389
rect 338 20355 422 20389
rect 237 20321 422 20355
rect 237 20287 304 20321
rect 338 20287 422 20321
rect 237 20253 422 20287
rect 237 20219 304 20253
rect 338 20219 422 20253
rect 237 20185 422 20219
rect 237 20151 304 20185
rect 338 20151 422 20185
rect 237 20117 422 20151
rect 237 20083 304 20117
rect 338 20083 422 20117
rect 237 20049 422 20083
rect 237 20015 304 20049
rect 338 20015 422 20049
rect 237 19981 422 20015
rect 237 19947 304 19981
rect 338 19947 422 19981
rect 237 19913 422 19947
rect 237 19879 304 19913
rect 338 19879 422 19913
rect 237 19845 422 19879
rect 237 19811 304 19845
rect 338 19811 422 19845
rect 237 19777 422 19811
rect 237 19743 304 19777
rect 338 19743 422 19777
rect 237 19709 422 19743
rect 237 19675 304 19709
rect 338 19675 422 19709
rect 237 19641 422 19675
rect 237 19607 304 19641
rect 338 19607 422 19641
rect 237 19573 422 19607
rect 237 19539 304 19573
rect 338 19539 422 19573
rect 237 19505 422 19539
rect 237 19471 304 19505
rect 338 19471 422 19505
rect 237 19437 422 19471
rect 237 19403 304 19437
rect 338 19403 422 19437
rect 237 19369 422 19403
rect 237 19335 304 19369
rect 338 19335 422 19369
rect 237 19301 422 19335
rect 237 19267 304 19301
rect 338 19267 422 19301
rect 237 19233 422 19267
rect 237 19199 304 19233
rect 338 19199 422 19233
rect 237 19165 422 19199
rect 237 19131 304 19165
rect 338 19131 422 19165
rect 237 19097 422 19131
rect 237 19063 304 19097
rect 338 19063 422 19097
rect 237 19029 422 19063
rect 237 18995 304 19029
rect 338 18995 422 19029
rect 237 18961 422 18995
rect 237 18927 304 18961
rect 338 18927 422 18961
rect 237 18893 422 18927
rect 237 18859 304 18893
rect 338 18859 422 18893
rect 237 18825 422 18859
rect 237 18791 304 18825
rect 338 18791 422 18825
rect 237 18757 422 18791
rect 237 18723 304 18757
rect 338 18723 422 18757
rect 237 18689 422 18723
rect 237 18655 304 18689
rect 338 18655 422 18689
rect 237 18621 422 18655
rect 237 18587 304 18621
rect 338 18587 422 18621
rect 237 18553 422 18587
rect 237 18519 304 18553
rect 338 18519 422 18553
rect 237 18485 422 18519
rect 237 18451 304 18485
rect 338 18451 422 18485
rect 237 18417 422 18451
rect 237 18383 304 18417
rect 338 18383 422 18417
rect 237 18349 422 18383
rect 237 18315 304 18349
rect 338 18315 422 18349
rect 237 18281 422 18315
rect 237 18247 304 18281
rect 338 18247 422 18281
rect 237 18213 422 18247
rect 237 18179 304 18213
rect 338 18179 422 18213
rect 237 18145 422 18179
rect 237 18111 304 18145
rect 338 18111 422 18145
rect 237 18077 422 18111
rect 237 18043 304 18077
rect 338 18043 422 18077
rect 237 18009 422 18043
rect 237 17975 304 18009
rect 338 17975 422 18009
rect 237 17941 422 17975
rect 237 17907 304 17941
rect 338 17907 422 17941
rect 237 17873 422 17907
rect 237 17839 304 17873
rect 338 17839 422 17873
rect 237 17805 422 17839
rect 237 17771 304 17805
rect 338 17771 422 17805
rect 237 17737 422 17771
rect 237 17703 304 17737
rect 338 17703 422 17737
rect 237 17669 422 17703
rect 237 17635 304 17669
rect 338 17635 422 17669
rect 237 17601 422 17635
rect 237 17567 304 17601
rect 338 17567 422 17601
rect 237 17533 422 17567
rect 237 17499 304 17533
rect 338 17499 422 17533
rect 237 17465 422 17499
rect 237 17431 304 17465
rect 338 17431 422 17465
rect 237 17397 422 17431
rect 237 17363 304 17397
rect 338 17363 422 17397
rect 237 17329 422 17363
rect 237 17295 304 17329
rect 338 17295 422 17329
rect 237 17261 422 17295
rect 237 17227 304 17261
rect 338 17227 422 17261
rect 237 17193 422 17227
rect 237 17159 304 17193
rect 338 17159 422 17193
rect 237 17125 422 17159
rect 237 17091 304 17125
rect 338 17091 422 17125
rect 237 17057 422 17091
rect 237 17023 304 17057
rect 338 17023 422 17057
rect 237 16989 422 17023
rect 237 16955 304 16989
rect 338 16955 422 16989
rect 237 16921 422 16955
rect 237 16887 304 16921
rect 338 16887 422 16921
rect 237 16853 422 16887
rect 237 16819 304 16853
rect 338 16819 422 16853
rect 237 16785 422 16819
rect 237 16751 304 16785
rect 338 16751 422 16785
rect 237 16717 422 16751
rect 237 16683 304 16717
rect 338 16683 422 16717
rect 237 16649 422 16683
rect 237 16615 304 16649
rect 338 16615 422 16649
rect 237 16581 422 16615
rect 237 16547 304 16581
rect 338 16547 422 16581
rect 237 16513 422 16547
rect 237 16479 304 16513
rect 338 16479 422 16513
rect 237 16445 422 16479
rect 237 16411 304 16445
rect 338 16411 422 16445
rect 237 16377 422 16411
rect 237 16343 304 16377
rect 338 16343 422 16377
rect 237 16309 422 16343
rect 237 16275 304 16309
rect 338 16275 422 16309
rect 237 16241 422 16275
rect 237 16207 304 16241
rect 338 16207 422 16241
rect 237 16173 422 16207
rect 237 16139 304 16173
rect 338 16139 422 16173
rect 237 16105 422 16139
rect 237 16071 304 16105
rect 338 16071 422 16105
rect 237 16037 422 16071
rect 237 16003 304 16037
rect 338 16003 422 16037
rect 237 15969 422 16003
rect 237 15935 304 15969
rect 338 15935 422 15969
rect 237 15901 422 15935
rect 237 15867 304 15901
rect 338 15867 422 15901
rect 237 15833 422 15867
rect 237 15799 304 15833
rect 338 15799 422 15833
rect 237 15765 422 15799
rect 237 15731 304 15765
rect 338 15731 422 15765
rect 237 15697 422 15731
rect 237 15663 304 15697
rect 338 15663 422 15697
rect 237 15629 422 15663
rect 237 15595 304 15629
rect 338 15595 422 15629
rect 237 15561 422 15595
rect 237 15527 304 15561
rect 338 15527 422 15561
rect 237 15493 422 15527
rect 237 15459 304 15493
rect 338 15459 422 15493
rect 237 15425 422 15459
rect 237 15391 304 15425
rect 338 15391 422 15425
rect 237 15357 422 15391
rect 237 15323 304 15357
rect 338 15323 422 15357
rect 237 15289 422 15323
rect 237 15255 304 15289
rect 338 15255 422 15289
rect 237 15221 422 15255
rect 237 15187 304 15221
rect 338 15187 422 15221
rect 237 15153 422 15187
rect 237 15119 304 15153
rect 338 15119 422 15153
rect 237 15085 422 15119
rect 237 15051 304 15085
rect 338 15051 422 15085
rect 237 15017 422 15051
rect 237 14983 304 15017
rect 338 14983 422 15017
rect 237 14949 422 14983
rect 237 14915 304 14949
rect 338 14915 422 14949
rect 237 14881 422 14915
rect 237 14847 304 14881
rect 338 14847 422 14881
rect 237 14813 422 14847
rect 237 14779 304 14813
rect 338 14779 422 14813
rect 237 14745 422 14779
rect 237 14711 304 14745
rect 338 14711 422 14745
rect 237 14677 422 14711
rect 1111 34692 13879 34734
rect 1111 34658 1297 34692
rect 1331 34658 1365 34692
rect 1399 34658 1433 34692
rect 1467 34658 1501 34692
rect 1535 34658 1569 34692
rect 1603 34658 1637 34692
rect 1671 34658 1705 34692
rect 1739 34658 1773 34692
rect 1807 34658 1841 34692
rect 1875 34658 1909 34692
rect 1943 34658 1977 34692
rect 2011 34658 2045 34692
rect 2079 34658 2113 34692
rect 2147 34658 2181 34692
rect 2215 34658 2249 34692
rect 2283 34658 2317 34692
rect 2351 34658 2385 34692
rect 2419 34658 2453 34692
rect 2487 34658 2521 34692
rect 2555 34658 2589 34692
rect 2623 34658 2657 34692
rect 2691 34658 2725 34692
rect 2759 34658 2793 34692
rect 2827 34658 2861 34692
rect 2895 34658 2929 34692
rect 2963 34658 2997 34692
rect 3031 34658 3065 34692
rect 3099 34658 3133 34692
rect 3167 34658 3201 34692
rect 3235 34658 3269 34692
rect 3303 34658 3337 34692
rect 3371 34658 3405 34692
rect 3439 34658 3473 34692
rect 3507 34658 3541 34692
rect 3575 34658 3609 34692
rect 3643 34658 3677 34692
rect 3711 34658 3745 34692
rect 3779 34658 3813 34692
rect 3847 34658 3881 34692
rect 3915 34658 3949 34692
rect 3983 34658 4017 34692
rect 4051 34658 4085 34692
rect 4119 34658 4153 34692
rect 4187 34658 4221 34692
rect 4255 34658 4289 34692
rect 4323 34658 4357 34692
rect 4391 34658 4425 34692
rect 4459 34658 4493 34692
rect 4527 34658 4561 34692
rect 4595 34658 4629 34692
rect 4663 34658 4697 34692
rect 4731 34658 4765 34692
rect 4799 34658 4833 34692
rect 4867 34658 4901 34692
rect 4935 34658 4969 34692
rect 5003 34658 5037 34692
rect 5071 34658 5105 34692
rect 5139 34658 5173 34692
rect 5207 34658 5241 34692
rect 5275 34658 5309 34692
rect 5343 34658 5377 34692
rect 5411 34658 5445 34692
rect 5479 34658 5513 34692
rect 5547 34658 5581 34692
rect 5615 34658 5649 34692
rect 5683 34658 5717 34692
rect 5751 34658 5785 34692
rect 5819 34658 5853 34692
rect 5887 34658 5921 34692
rect 5955 34658 5989 34692
rect 6023 34658 6057 34692
rect 6091 34658 6125 34692
rect 6159 34658 6193 34692
rect 6227 34658 6261 34692
rect 6295 34658 6329 34692
rect 6363 34658 6397 34692
rect 6431 34658 6465 34692
rect 6499 34658 6533 34692
rect 6567 34658 6601 34692
rect 6635 34658 6669 34692
rect 6703 34658 6737 34692
rect 6771 34658 6805 34692
rect 6839 34658 6873 34692
rect 6907 34658 6941 34692
rect 6975 34658 7009 34692
rect 7043 34658 7077 34692
rect 7111 34658 7145 34692
rect 7179 34658 7213 34692
rect 7247 34658 7281 34692
rect 7315 34658 7349 34692
rect 7383 34658 7417 34692
rect 7451 34658 7485 34692
rect 7519 34658 7553 34692
rect 7587 34658 7621 34692
rect 7655 34658 7689 34692
rect 7723 34658 7757 34692
rect 7791 34658 7825 34692
rect 7859 34658 7893 34692
rect 7927 34658 7961 34692
rect 7995 34658 8029 34692
rect 8063 34658 8097 34692
rect 8131 34658 8165 34692
rect 8199 34658 8233 34692
rect 8267 34658 8301 34692
rect 8335 34658 8369 34692
rect 8403 34658 8437 34692
rect 8471 34658 8505 34692
rect 8539 34658 8573 34692
rect 8607 34658 8641 34692
rect 8675 34658 8709 34692
rect 8743 34658 8777 34692
rect 8811 34658 8845 34692
rect 8879 34658 8913 34692
rect 8947 34658 8981 34692
rect 9015 34658 9049 34692
rect 9083 34658 9117 34692
rect 9151 34658 9185 34692
rect 9219 34658 9253 34692
rect 9287 34658 9321 34692
rect 9355 34658 9389 34692
rect 9423 34658 9457 34692
rect 9491 34658 9525 34692
rect 9559 34658 9593 34692
rect 9627 34658 9661 34692
rect 9695 34658 9729 34692
rect 9763 34658 9797 34692
rect 9831 34658 9865 34692
rect 9899 34658 9933 34692
rect 9967 34658 10001 34692
rect 10035 34658 10069 34692
rect 10103 34658 10137 34692
rect 10171 34658 10205 34692
rect 10239 34658 10273 34692
rect 10307 34658 10341 34692
rect 10375 34658 10409 34692
rect 10443 34658 10477 34692
rect 10511 34658 10545 34692
rect 10579 34658 10613 34692
rect 10647 34658 10681 34692
rect 10715 34658 10749 34692
rect 10783 34658 10817 34692
rect 10851 34658 10885 34692
rect 10919 34658 10953 34692
rect 10987 34658 11021 34692
rect 11055 34658 11089 34692
rect 11123 34658 11157 34692
rect 11191 34658 11225 34692
rect 11259 34658 11293 34692
rect 11327 34658 11361 34692
rect 11395 34658 11429 34692
rect 11463 34658 11497 34692
rect 11531 34658 11565 34692
rect 11599 34658 11633 34692
rect 11667 34658 11701 34692
rect 11735 34658 11769 34692
rect 11803 34658 11837 34692
rect 11871 34658 11905 34692
rect 11939 34658 11973 34692
rect 12007 34658 12041 34692
rect 12075 34658 12109 34692
rect 12143 34658 12177 34692
rect 12211 34658 12245 34692
rect 12279 34658 12313 34692
rect 12347 34658 12381 34692
rect 12415 34658 12449 34692
rect 12483 34658 12517 34692
rect 12551 34658 12585 34692
rect 12619 34658 12653 34692
rect 12687 34658 12721 34692
rect 12755 34658 12789 34692
rect 12823 34658 12857 34692
rect 12891 34658 12925 34692
rect 12959 34658 12993 34692
rect 13027 34658 13061 34692
rect 13095 34658 13129 34692
rect 13163 34658 13197 34692
rect 13231 34658 13265 34692
rect 13299 34658 13333 34692
rect 13367 34658 13401 34692
rect 13435 34658 13469 34692
rect 13503 34658 13537 34692
rect 13571 34658 13605 34692
rect 13639 34658 13673 34692
rect 13707 34658 13879 34692
rect 1111 34616 13879 34658
rect 1111 34475 1229 34616
rect 1111 34441 1153 34475
rect 1187 34441 1229 34475
rect 1111 34407 1229 34441
rect 1111 34373 1153 34407
rect 1187 34373 1229 34407
rect 1111 34339 1229 34373
rect 1111 34305 1153 34339
rect 1187 34305 1229 34339
rect 1111 34271 1229 34305
rect 1111 34237 1153 34271
rect 1187 34237 1229 34271
rect 1111 34203 1229 34237
rect 1111 34169 1153 34203
rect 1187 34169 1229 34203
rect 1111 34135 1229 34169
rect 1111 34101 1153 34135
rect 1187 34101 1229 34135
rect 1111 34067 1229 34101
rect 1111 34033 1153 34067
rect 1187 34033 1229 34067
rect 1111 33999 1229 34033
rect 1111 33965 1153 33999
rect 1187 33965 1229 33999
rect 1111 33931 1229 33965
rect 1111 33897 1153 33931
rect 1187 33897 1229 33931
rect 1111 33863 1229 33897
rect 1111 33829 1153 33863
rect 1187 33829 1229 33863
rect 1111 33795 1229 33829
rect 1111 33761 1153 33795
rect 1187 33761 1229 33795
rect 1111 33727 1229 33761
rect 1111 33693 1153 33727
rect 1187 33693 1229 33727
rect 1111 33659 1229 33693
rect 1111 33625 1153 33659
rect 1187 33625 1229 33659
rect 1111 33591 1229 33625
rect 1111 33557 1153 33591
rect 1187 33557 1229 33591
rect 1111 33523 1229 33557
rect 1111 33489 1153 33523
rect 1187 33489 1229 33523
rect 1111 33455 1229 33489
rect 1111 33421 1153 33455
rect 1187 33421 1229 33455
rect 1111 33387 1229 33421
rect 1111 33353 1153 33387
rect 1187 33353 1229 33387
rect 1111 33319 1229 33353
rect 1111 33285 1153 33319
rect 1187 33285 1229 33319
rect 1111 33251 1229 33285
rect 1111 33217 1153 33251
rect 1187 33217 1229 33251
rect 1111 33183 1229 33217
rect 1111 33149 1153 33183
rect 1187 33149 1229 33183
rect 1111 33115 1229 33149
rect 1111 33081 1153 33115
rect 1187 33081 1229 33115
rect 1111 33047 1229 33081
rect 1111 33013 1153 33047
rect 1187 33013 1229 33047
rect 1111 32979 1229 33013
rect 1111 32945 1153 32979
rect 1187 32945 1229 32979
rect 1111 32911 1229 32945
rect 1111 32877 1153 32911
rect 1187 32877 1229 32911
rect 1111 32843 1229 32877
rect 1111 32809 1153 32843
rect 1187 32809 1229 32843
rect 1111 32775 1229 32809
rect 1111 32741 1153 32775
rect 1187 32741 1229 32775
rect 1111 32707 1229 32741
rect 1111 32673 1153 32707
rect 1187 32673 1229 32707
rect 1111 32639 1229 32673
rect 1111 32605 1153 32639
rect 1187 32605 1229 32639
rect 1111 32571 1229 32605
rect 1111 32537 1153 32571
rect 1187 32537 1229 32571
rect 1111 32503 1229 32537
rect 1111 32469 1153 32503
rect 1187 32469 1229 32503
rect 1111 32435 1229 32469
rect 1111 32401 1153 32435
rect 1187 32401 1229 32435
rect 1111 32367 1229 32401
rect 1111 32333 1153 32367
rect 1187 32333 1229 32367
rect 1111 32299 1229 32333
rect 1111 32265 1153 32299
rect 1187 32265 1229 32299
rect 1111 32231 1229 32265
rect 1111 32197 1153 32231
rect 1187 32197 1229 32231
rect 1111 32163 1229 32197
rect 1111 32129 1153 32163
rect 1187 32129 1229 32163
rect 1111 32095 1229 32129
rect 1111 32061 1153 32095
rect 1187 32061 1229 32095
rect 1111 32027 1229 32061
rect 1111 31993 1153 32027
rect 1187 31993 1229 32027
rect 1111 31959 1229 31993
rect 1111 31925 1153 31959
rect 1187 31925 1229 31959
rect 1111 31891 1229 31925
rect 1111 31857 1153 31891
rect 1187 31857 1229 31891
rect 1111 31823 1229 31857
rect 1111 31789 1153 31823
rect 1187 31789 1229 31823
rect 1111 31755 1229 31789
rect 1111 31721 1153 31755
rect 1187 31721 1229 31755
rect 1111 31687 1229 31721
rect 1111 31653 1153 31687
rect 1187 31653 1229 31687
rect 1111 31619 1229 31653
rect 1111 31585 1153 31619
rect 1187 31585 1229 31619
rect 1111 31551 1229 31585
rect 1111 31517 1153 31551
rect 1187 31517 1229 31551
rect 1111 31483 1229 31517
rect 1111 31449 1153 31483
rect 1187 31449 1229 31483
rect 1111 31415 1229 31449
rect 1111 31381 1153 31415
rect 1187 31381 1229 31415
rect 1111 31347 1229 31381
rect 1111 31313 1153 31347
rect 1187 31313 1229 31347
rect 1111 31279 1229 31313
rect 1111 31245 1153 31279
rect 1187 31245 1229 31279
rect 1111 31211 1229 31245
rect 1111 31177 1153 31211
rect 1187 31177 1229 31211
rect 1111 31143 1229 31177
rect 1111 31109 1153 31143
rect 1187 31109 1229 31143
rect 1111 31075 1229 31109
rect 1111 31041 1153 31075
rect 1187 31041 1229 31075
rect 1111 31007 1229 31041
rect 1111 30973 1153 31007
rect 1187 30973 1229 31007
rect 1111 30939 1229 30973
rect 1111 30905 1153 30939
rect 1187 30905 1229 30939
rect 1111 30871 1229 30905
rect 1111 30837 1153 30871
rect 1187 30837 1229 30871
rect 1111 30803 1229 30837
rect 1111 30769 1153 30803
rect 1187 30769 1229 30803
rect 1111 30735 1229 30769
rect 1111 30701 1153 30735
rect 1187 30701 1229 30735
rect 1111 30667 1229 30701
rect 1111 30633 1153 30667
rect 1187 30633 1229 30667
rect 1111 30599 1229 30633
rect 1111 30565 1153 30599
rect 1187 30565 1229 30599
rect 1111 30531 1229 30565
rect 1111 30497 1153 30531
rect 1187 30497 1229 30531
rect 1111 30463 1229 30497
rect 1111 30429 1153 30463
rect 1187 30429 1229 30463
rect 1111 30395 1229 30429
rect 1111 30361 1153 30395
rect 1187 30361 1229 30395
rect 1111 30327 1229 30361
rect 1111 30293 1153 30327
rect 1187 30293 1229 30327
rect 1111 30259 1229 30293
rect 1111 30225 1153 30259
rect 1187 30225 1229 30259
rect 1111 30191 1229 30225
rect 1111 30157 1153 30191
rect 1187 30157 1229 30191
rect 1111 30123 1229 30157
rect 1111 30089 1153 30123
rect 1187 30089 1229 30123
rect 1111 30055 1229 30089
rect 1111 30021 1153 30055
rect 1187 30021 1229 30055
rect 1111 29987 1229 30021
rect 1111 29953 1153 29987
rect 1187 29953 1229 29987
rect 1111 29919 1229 29953
rect 1111 29885 1153 29919
rect 1187 29885 1229 29919
rect 1111 29851 1229 29885
rect 1111 29817 1153 29851
rect 1187 29817 1229 29851
rect 1111 29783 1229 29817
rect 1111 29749 1153 29783
rect 1187 29749 1229 29783
rect 1111 29715 1229 29749
rect 1111 29681 1153 29715
rect 1187 29681 1229 29715
rect 1111 29647 1229 29681
rect 1111 29613 1153 29647
rect 1187 29613 1229 29647
rect 1111 29579 1229 29613
rect 1111 29545 1153 29579
rect 1187 29545 1229 29579
rect 1111 29511 1229 29545
rect 1111 29477 1153 29511
rect 1187 29477 1229 29511
rect 1111 29443 1229 29477
rect 1111 29409 1153 29443
rect 1187 29409 1229 29443
rect 1111 29375 1229 29409
rect 1111 29341 1153 29375
rect 1187 29341 1229 29375
rect 1111 29307 1229 29341
rect 1111 29273 1153 29307
rect 1187 29273 1229 29307
rect 1111 29239 1229 29273
rect 1111 29205 1153 29239
rect 1187 29205 1229 29239
rect 1111 29171 1229 29205
rect 1111 29137 1153 29171
rect 1187 29137 1229 29171
rect 1111 29103 1229 29137
rect 1111 29069 1153 29103
rect 1187 29069 1229 29103
rect 1111 29035 1229 29069
rect 1111 29001 1153 29035
rect 1187 29001 1229 29035
rect 1111 28967 1229 29001
rect 1111 28933 1153 28967
rect 1187 28933 1229 28967
rect 1111 28899 1229 28933
rect 13761 34470 13879 34616
rect 13761 34436 13801 34470
rect 13835 34436 13879 34470
rect 13761 34402 13879 34436
rect 13761 34368 13801 34402
rect 13835 34368 13879 34402
rect 13761 34334 13879 34368
rect 13761 34300 13801 34334
rect 13835 34300 13879 34334
rect 13761 34266 13879 34300
rect 13761 34232 13801 34266
rect 13835 34232 13879 34266
rect 13761 34198 13879 34232
rect 13761 34164 13801 34198
rect 13835 34164 13879 34198
rect 13761 34130 13879 34164
rect 13761 34096 13801 34130
rect 13835 34096 13879 34130
rect 13761 34062 13879 34096
rect 13761 34028 13801 34062
rect 13835 34028 13879 34062
rect 13761 33994 13879 34028
rect 13761 33960 13801 33994
rect 13835 33960 13879 33994
rect 13761 33926 13879 33960
rect 13761 33892 13801 33926
rect 13835 33892 13879 33926
rect 13761 33858 13879 33892
rect 13761 33824 13801 33858
rect 13835 33824 13879 33858
rect 13761 33790 13879 33824
rect 13761 33756 13801 33790
rect 13835 33756 13879 33790
rect 13761 33722 13879 33756
rect 13761 33688 13801 33722
rect 13835 33688 13879 33722
rect 13761 33654 13879 33688
rect 13761 33620 13801 33654
rect 13835 33620 13879 33654
rect 13761 33586 13879 33620
rect 13761 33552 13801 33586
rect 13835 33552 13879 33586
rect 13761 33518 13879 33552
rect 13761 33484 13801 33518
rect 13835 33484 13879 33518
rect 13761 33450 13879 33484
rect 13761 33416 13801 33450
rect 13835 33416 13879 33450
rect 13761 33382 13879 33416
rect 13761 33348 13801 33382
rect 13835 33348 13879 33382
rect 13761 33314 13879 33348
rect 13761 33280 13801 33314
rect 13835 33280 13879 33314
rect 13761 33246 13879 33280
rect 13761 33212 13801 33246
rect 13835 33212 13879 33246
rect 13761 33178 13879 33212
rect 13761 33144 13801 33178
rect 13835 33144 13879 33178
rect 13761 33110 13879 33144
rect 13761 33076 13801 33110
rect 13835 33076 13879 33110
rect 13761 33042 13879 33076
rect 13761 33008 13801 33042
rect 13835 33008 13879 33042
rect 13761 32974 13879 33008
rect 13761 32940 13801 32974
rect 13835 32940 13879 32974
rect 13761 32906 13879 32940
rect 13761 32872 13801 32906
rect 13835 32872 13879 32906
rect 13761 32838 13879 32872
rect 13761 32804 13801 32838
rect 13835 32804 13879 32838
rect 13761 32770 13879 32804
rect 13761 32736 13801 32770
rect 13835 32736 13879 32770
rect 13761 32702 13879 32736
rect 13761 32668 13801 32702
rect 13835 32668 13879 32702
rect 13761 32634 13879 32668
rect 13761 32600 13801 32634
rect 13835 32600 13879 32634
rect 13761 32566 13879 32600
rect 13761 32532 13801 32566
rect 13835 32532 13879 32566
rect 13761 32498 13879 32532
rect 13761 32464 13801 32498
rect 13835 32464 13879 32498
rect 13761 32430 13879 32464
rect 13761 32396 13801 32430
rect 13835 32396 13879 32430
rect 13761 32362 13879 32396
rect 13761 32328 13801 32362
rect 13835 32328 13879 32362
rect 13761 32294 13879 32328
rect 13761 32260 13801 32294
rect 13835 32260 13879 32294
rect 13761 32226 13879 32260
rect 13761 32192 13801 32226
rect 13835 32192 13879 32226
rect 13761 32158 13879 32192
rect 13761 32124 13801 32158
rect 13835 32124 13879 32158
rect 13761 32090 13879 32124
rect 13761 32056 13801 32090
rect 13835 32056 13879 32090
rect 13761 32022 13879 32056
rect 13761 31988 13801 32022
rect 13835 31988 13879 32022
rect 13761 31954 13879 31988
rect 13761 31920 13801 31954
rect 13835 31920 13879 31954
rect 13761 31886 13879 31920
rect 13761 31852 13801 31886
rect 13835 31852 13879 31886
rect 13761 31818 13879 31852
rect 13761 31784 13801 31818
rect 13835 31784 13879 31818
rect 13761 31750 13879 31784
rect 13761 31716 13801 31750
rect 13835 31716 13879 31750
rect 13761 31682 13879 31716
rect 13761 31648 13801 31682
rect 13835 31648 13879 31682
rect 13761 31614 13879 31648
rect 13761 31580 13801 31614
rect 13835 31580 13879 31614
rect 13761 31546 13879 31580
rect 13761 31512 13801 31546
rect 13835 31512 13879 31546
rect 13761 31478 13879 31512
rect 13761 31444 13801 31478
rect 13835 31444 13879 31478
rect 13761 31410 13879 31444
rect 13761 31376 13801 31410
rect 13835 31376 13879 31410
rect 13761 31342 13879 31376
rect 13761 31308 13801 31342
rect 13835 31308 13879 31342
rect 13761 31274 13879 31308
rect 13761 31240 13801 31274
rect 13835 31240 13879 31274
rect 13761 31206 13879 31240
rect 13761 31172 13801 31206
rect 13835 31172 13879 31206
rect 13761 31138 13879 31172
rect 13761 31104 13801 31138
rect 13835 31104 13879 31138
rect 13761 31070 13879 31104
rect 13761 31036 13801 31070
rect 13835 31036 13879 31070
rect 13761 31002 13879 31036
rect 13761 30968 13801 31002
rect 13835 30968 13879 31002
rect 13761 30934 13879 30968
rect 13761 30900 13801 30934
rect 13835 30900 13879 30934
rect 13761 30866 13879 30900
rect 13761 30832 13801 30866
rect 13835 30832 13879 30866
rect 13761 30798 13879 30832
rect 13761 30764 13801 30798
rect 13835 30764 13879 30798
rect 13761 30730 13879 30764
rect 13761 30696 13801 30730
rect 13835 30696 13879 30730
rect 13761 30662 13879 30696
rect 13761 30628 13801 30662
rect 13835 30628 13879 30662
rect 13761 30594 13879 30628
rect 13761 30560 13801 30594
rect 13835 30560 13879 30594
rect 13761 30526 13879 30560
rect 13761 30492 13801 30526
rect 13835 30492 13879 30526
rect 13761 30458 13879 30492
rect 13761 30424 13801 30458
rect 13835 30424 13879 30458
rect 13761 30390 13879 30424
rect 13761 30356 13801 30390
rect 13835 30356 13879 30390
rect 13761 30322 13879 30356
rect 13761 30288 13801 30322
rect 13835 30288 13879 30322
rect 13761 30254 13879 30288
rect 13761 30220 13801 30254
rect 13835 30220 13879 30254
rect 13761 30186 13879 30220
rect 13761 30152 13801 30186
rect 13835 30152 13879 30186
rect 13761 30118 13879 30152
rect 13761 30084 13801 30118
rect 13835 30084 13879 30118
rect 13761 30050 13879 30084
rect 13761 30016 13801 30050
rect 13835 30016 13879 30050
rect 13761 29982 13879 30016
rect 13761 29948 13801 29982
rect 13835 29948 13879 29982
rect 13761 29914 13879 29948
rect 13761 29880 13801 29914
rect 13835 29880 13879 29914
rect 13761 29846 13879 29880
rect 13761 29812 13801 29846
rect 13835 29812 13879 29846
rect 13761 29778 13879 29812
rect 13761 29744 13801 29778
rect 13835 29744 13879 29778
rect 13761 29710 13879 29744
rect 13761 29676 13801 29710
rect 13835 29676 13879 29710
rect 13761 29642 13879 29676
rect 13761 29608 13801 29642
rect 13835 29608 13879 29642
rect 13761 29574 13879 29608
rect 13761 29540 13801 29574
rect 13835 29540 13879 29574
rect 13761 29506 13879 29540
rect 13761 29472 13801 29506
rect 13835 29472 13879 29506
rect 13761 29438 13879 29472
rect 13761 29404 13801 29438
rect 13835 29404 13879 29438
rect 13761 29370 13879 29404
rect 13761 29336 13801 29370
rect 13835 29336 13879 29370
rect 13761 29302 13879 29336
rect 13761 29268 13801 29302
rect 13835 29268 13879 29302
rect 13761 29234 13879 29268
rect 13761 29200 13801 29234
rect 13835 29200 13879 29234
rect 13761 29166 13879 29200
rect 13761 29132 13801 29166
rect 13835 29132 13879 29166
rect 13761 29098 13879 29132
rect 13761 29064 13801 29098
rect 13835 29064 13879 29098
rect 13761 29030 13879 29064
rect 13761 28996 13801 29030
rect 13835 28996 13879 29030
rect 13761 28962 13879 28996
rect 13761 28928 13801 28962
rect 13835 28928 13879 28962
rect 1111 28865 1153 28899
rect 1187 28865 1229 28899
rect 1111 28831 1229 28865
rect 1111 28797 1153 28831
rect 1187 28797 1229 28831
rect 1111 28763 1229 28797
rect 1111 28729 1153 28763
rect 1187 28729 1229 28763
rect 1111 28695 1229 28729
rect 1111 28661 1153 28695
rect 1187 28661 1229 28695
rect 1111 28627 1229 28661
rect 1111 28593 1153 28627
rect 1187 28593 1229 28627
rect 1111 28559 1229 28593
rect 1111 28525 1153 28559
rect 1187 28525 1229 28559
rect 1111 28491 1229 28525
rect 1111 28457 1153 28491
rect 1187 28457 1229 28491
rect 1111 28423 1229 28457
rect 1111 28389 1153 28423
rect 1187 28389 1229 28423
rect 1111 28355 1229 28389
rect 1111 28321 1153 28355
rect 1187 28321 1229 28355
rect 1111 28287 1229 28321
rect 1111 28253 1153 28287
rect 1187 28253 1229 28287
rect 1111 28219 1229 28253
rect 1111 28185 1153 28219
rect 1187 28185 1229 28219
rect 1111 28151 1229 28185
rect 1111 28117 1153 28151
rect 1187 28117 1229 28151
rect 1111 28083 1229 28117
rect 1111 28049 1153 28083
rect 1187 28049 1229 28083
rect 1111 28015 1229 28049
rect 1111 27981 1153 28015
rect 1187 27981 1229 28015
rect 1111 27947 1229 27981
rect 1111 27913 1153 27947
rect 1187 27913 1229 27947
rect 1111 27879 1229 27913
rect 1111 27845 1153 27879
rect 1187 27845 1229 27879
rect 1111 27811 1229 27845
rect 1111 27777 1153 27811
rect 1187 27777 1229 27811
rect 1111 27743 1229 27777
rect 1111 27709 1153 27743
rect 1187 27709 1229 27743
rect 1111 27675 1229 27709
rect 1111 27641 1153 27675
rect 1187 27641 1229 27675
rect 1111 27607 1229 27641
rect 1111 27573 1153 27607
rect 1187 27573 1229 27607
rect 1111 27539 1229 27573
rect 1111 27505 1153 27539
rect 1187 27505 1229 27539
rect 1111 27471 1229 27505
rect 1111 27437 1153 27471
rect 1187 27437 1229 27471
rect 1111 27403 1229 27437
rect 1111 27369 1153 27403
rect 1187 27369 1229 27403
rect 1111 27335 1229 27369
rect 1111 27301 1153 27335
rect 1187 27301 1229 27335
rect 1111 27267 1229 27301
rect 1111 27233 1153 27267
rect 1187 27233 1229 27267
rect 1111 27199 1229 27233
rect 1111 27165 1153 27199
rect 1187 27165 1229 27199
rect 1111 27131 1229 27165
rect 1111 27097 1153 27131
rect 1187 27097 1229 27131
rect 1111 27063 1229 27097
rect 1111 27029 1153 27063
rect 1187 27029 1229 27063
rect 2364 28273 12636 28289
rect 2364 28239 2485 28273
rect 2519 28239 2553 28273
rect 2587 28239 2621 28273
rect 2655 28239 2689 28273
rect 2723 28239 2757 28273
rect 2791 28239 2825 28273
rect 2859 28239 2893 28273
rect 2927 28239 2961 28273
rect 2995 28239 3029 28273
rect 3063 28239 3097 28273
rect 3131 28239 3165 28273
rect 3199 28239 3233 28273
rect 3267 28239 3301 28273
rect 3335 28239 3369 28273
rect 3403 28239 3437 28273
rect 3471 28239 3505 28273
rect 3539 28239 3573 28273
rect 3607 28239 3641 28273
rect 3675 28239 3709 28273
rect 3743 28239 3777 28273
rect 3811 28239 3845 28273
rect 3879 28239 3913 28273
rect 3947 28239 3981 28273
rect 4015 28239 4049 28273
rect 4083 28239 4117 28273
rect 4151 28239 4185 28273
rect 4219 28239 4253 28273
rect 4287 28239 4321 28273
rect 4355 28239 4389 28273
rect 4423 28239 4457 28273
rect 4491 28239 4525 28273
rect 4559 28239 4593 28273
rect 4627 28239 4661 28273
rect 4695 28239 4729 28273
rect 4763 28239 4797 28273
rect 4831 28239 4865 28273
rect 4899 28239 4933 28273
rect 4967 28239 5001 28273
rect 5035 28239 5069 28273
rect 5103 28239 5137 28273
rect 5171 28239 5205 28273
rect 5239 28239 5273 28273
rect 5307 28239 5341 28273
rect 5375 28239 5409 28273
rect 5443 28239 5477 28273
rect 5511 28239 5545 28273
rect 5579 28239 5613 28273
rect 5647 28239 5681 28273
rect 5715 28239 5749 28273
rect 5783 28239 5817 28273
rect 5851 28239 5885 28273
rect 5919 28239 5953 28273
rect 5987 28239 6021 28273
rect 6055 28239 6089 28273
rect 6123 28239 6157 28273
rect 6191 28239 6225 28273
rect 6259 28239 6293 28273
rect 6327 28239 6361 28273
rect 6395 28239 6429 28273
rect 6463 28239 6497 28273
rect 6531 28239 6565 28273
rect 6599 28239 6633 28273
rect 6667 28239 6701 28273
rect 6735 28239 6769 28273
rect 6803 28239 6837 28273
rect 6871 28239 6905 28273
rect 6939 28239 6973 28273
rect 7007 28239 7041 28273
rect 7075 28239 7109 28273
rect 7143 28239 7177 28273
rect 7211 28239 7245 28273
rect 7279 28239 7313 28273
rect 7347 28239 7381 28273
rect 7415 28239 7449 28273
rect 7483 28239 7517 28273
rect 7551 28239 7585 28273
rect 7619 28239 7653 28273
rect 7687 28239 7721 28273
rect 7755 28239 7789 28273
rect 7823 28239 7857 28273
rect 7891 28239 7925 28273
rect 7959 28239 7993 28273
rect 8027 28239 8061 28273
rect 8095 28239 8129 28273
rect 8163 28239 8197 28273
rect 8231 28239 8265 28273
rect 8299 28239 8333 28273
rect 8367 28239 8401 28273
rect 8435 28239 8469 28273
rect 8503 28239 8537 28273
rect 8571 28239 8605 28273
rect 8639 28239 8673 28273
rect 8707 28239 8741 28273
rect 8775 28239 8809 28273
rect 8843 28239 8877 28273
rect 8911 28239 8945 28273
rect 8979 28239 9013 28273
rect 9047 28239 9081 28273
rect 9115 28239 9149 28273
rect 9183 28239 9217 28273
rect 9251 28239 9285 28273
rect 9319 28239 9353 28273
rect 9387 28239 9421 28273
rect 9455 28239 9489 28273
rect 9523 28239 9557 28273
rect 9591 28239 9625 28273
rect 9659 28239 9693 28273
rect 9727 28239 9761 28273
rect 9795 28239 9829 28273
rect 9863 28239 9897 28273
rect 9931 28239 9965 28273
rect 9999 28239 10033 28273
rect 10067 28239 10101 28273
rect 10135 28239 10169 28273
rect 10203 28239 10237 28273
rect 10271 28239 10305 28273
rect 10339 28239 10373 28273
rect 10407 28239 10441 28273
rect 10475 28239 10509 28273
rect 10543 28239 10577 28273
rect 10611 28239 10645 28273
rect 10679 28239 10713 28273
rect 10747 28239 10781 28273
rect 10815 28239 10849 28273
rect 10883 28239 10917 28273
rect 10951 28239 10985 28273
rect 11019 28239 11053 28273
rect 11087 28239 11121 28273
rect 11155 28239 11189 28273
rect 11223 28239 11257 28273
rect 11291 28239 11325 28273
rect 11359 28239 11393 28273
rect 11427 28239 11461 28273
rect 11495 28239 11529 28273
rect 11563 28239 11597 28273
rect 11631 28239 11665 28273
rect 11699 28239 11733 28273
rect 11767 28239 11801 28273
rect 11835 28239 11869 28273
rect 11903 28239 11937 28273
rect 11971 28239 12005 28273
rect 12039 28239 12073 28273
rect 12107 28239 12141 28273
rect 12175 28239 12209 28273
rect 12243 28239 12277 28273
rect 12311 28239 12345 28273
rect 12379 28239 12413 28273
rect 12447 28239 12481 28273
rect 12515 28239 12636 28273
rect 2364 28203 12636 28239
rect 2364 28169 2485 28203
rect 2519 28169 2553 28203
rect 2587 28169 2621 28203
rect 2655 28169 2689 28203
rect 2723 28169 2757 28203
rect 2791 28169 2825 28203
rect 2859 28169 2893 28203
rect 2927 28169 2961 28203
rect 2995 28169 3029 28203
rect 3063 28169 3097 28203
rect 3131 28169 3165 28203
rect 3199 28169 3233 28203
rect 3267 28169 3301 28203
rect 3335 28169 3369 28203
rect 3403 28169 3437 28203
rect 3471 28169 3505 28203
rect 3539 28169 3573 28203
rect 3607 28169 3641 28203
rect 3675 28169 3709 28203
rect 3743 28169 3777 28203
rect 3811 28169 3845 28203
rect 3879 28169 3913 28203
rect 3947 28169 3981 28203
rect 4015 28169 4049 28203
rect 4083 28169 4117 28203
rect 4151 28169 4185 28203
rect 4219 28169 4253 28203
rect 4287 28169 4321 28203
rect 4355 28169 4389 28203
rect 4423 28169 4457 28203
rect 4491 28169 4525 28203
rect 4559 28169 4593 28203
rect 4627 28169 4661 28203
rect 4695 28169 4729 28203
rect 4763 28169 4797 28203
rect 4831 28169 4865 28203
rect 4899 28169 4933 28203
rect 4967 28169 5001 28203
rect 5035 28169 5069 28203
rect 5103 28169 5137 28203
rect 5171 28169 5205 28203
rect 5239 28169 5273 28203
rect 5307 28169 5341 28203
rect 5375 28169 5409 28203
rect 5443 28169 5477 28203
rect 5511 28169 5545 28203
rect 5579 28169 5613 28203
rect 5647 28169 5681 28203
rect 5715 28169 5749 28203
rect 5783 28169 5817 28203
rect 5851 28169 5885 28203
rect 5919 28169 5953 28203
rect 5987 28169 6021 28203
rect 6055 28169 6089 28203
rect 6123 28169 6157 28203
rect 6191 28169 6225 28203
rect 6259 28169 6293 28203
rect 6327 28169 6361 28203
rect 6395 28169 6429 28203
rect 6463 28169 6497 28203
rect 6531 28169 6565 28203
rect 6599 28169 6633 28203
rect 6667 28169 6701 28203
rect 6735 28169 6769 28203
rect 6803 28169 6837 28203
rect 6871 28169 6905 28203
rect 6939 28169 6973 28203
rect 7007 28169 7041 28203
rect 7075 28169 7109 28203
rect 7143 28169 7177 28203
rect 7211 28169 7245 28203
rect 7279 28169 7313 28203
rect 7347 28169 7381 28203
rect 7415 28169 7449 28203
rect 7483 28169 7517 28203
rect 7551 28169 7585 28203
rect 7619 28169 7653 28203
rect 7687 28169 7721 28203
rect 7755 28169 7789 28203
rect 7823 28169 7857 28203
rect 7891 28169 7925 28203
rect 7959 28169 7993 28203
rect 8027 28169 8061 28203
rect 8095 28169 8129 28203
rect 8163 28169 8197 28203
rect 8231 28169 8265 28203
rect 8299 28169 8333 28203
rect 8367 28169 8401 28203
rect 8435 28169 8469 28203
rect 8503 28169 8537 28203
rect 8571 28169 8605 28203
rect 8639 28169 8673 28203
rect 8707 28169 8741 28203
rect 8775 28169 8809 28203
rect 8843 28169 8877 28203
rect 8911 28169 8945 28203
rect 8979 28169 9013 28203
rect 9047 28169 9081 28203
rect 9115 28169 9149 28203
rect 9183 28169 9217 28203
rect 9251 28169 9285 28203
rect 9319 28169 9353 28203
rect 9387 28169 9421 28203
rect 9455 28169 9489 28203
rect 9523 28169 9557 28203
rect 9591 28169 9625 28203
rect 9659 28169 9693 28203
rect 9727 28169 9761 28203
rect 9795 28169 9829 28203
rect 9863 28169 9897 28203
rect 9931 28169 9965 28203
rect 9999 28169 10033 28203
rect 10067 28169 10101 28203
rect 10135 28169 10169 28203
rect 10203 28169 10237 28203
rect 10271 28169 10305 28203
rect 10339 28169 10373 28203
rect 10407 28169 10441 28203
rect 10475 28169 10509 28203
rect 10543 28169 10577 28203
rect 10611 28169 10645 28203
rect 10679 28169 10713 28203
rect 10747 28169 10781 28203
rect 10815 28169 10849 28203
rect 10883 28169 10917 28203
rect 10951 28169 10985 28203
rect 11019 28169 11053 28203
rect 11087 28169 11121 28203
rect 11155 28169 11189 28203
rect 11223 28169 11257 28203
rect 11291 28169 11325 28203
rect 11359 28169 11393 28203
rect 11427 28169 11461 28203
rect 11495 28169 11529 28203
rect 11563 28169 11597 28203
rect 11631 28169 11665 28203
rect 11699 28169 11733 28203
rect 11767 28169 11801 28203
rect 11835 28169 11869 28203
rect 11903 28169 11937 28203
rect 11971 28169 12005 28203
rect 12039 28169 12073 28203
rect 12107 28169 12141 28203
rect 12175 28169 12209 28203
rect 12243 28169 12277 28203
rect 12311 28169 12345 28203
rect 12379 28169 12413 28203
rect 12447 28169 12481 28203
rect 12515 28169 12636 28203
rect 2364 28157 12636 28169
rect 2364 28098 2422 28157
rect 2364 28064 2376 28098
rect 2410 28064 2422 28098
rect 12578 28098 12636 28157
rect 2364 28030 2422 28064
rect 2364 27996 2376 28030
rect 2410 27996 2422 28030
rect 2364 27962 2422 27996
rect 2364 27928 2376 27962
rect 2410 27928 2422 27962
rect 2364 27894 2422 27928
rect 2364 27860 2376 27894
rect 2410 27860 2422 27894
rect 12578 28064 12590 28098
rect 12624 28064 12636 28098
rect 12578 28030 12636 28064
rect 12578 27996 12590 28030
rect 12624 27996 12636 28030
rect 12578 27962 12636 27996
rect 12578 27928 12590 27962
rect 12624 27928 12636 27962
rect 12578 27894 12636 27928
rect 2364 27801 2422 27860
rect 12578 27860 12590 27894
rect 12624 27860 12636 27894
rect 12578 27801 12636 27860
rect 2364 27789 12636 27801
rect 2364 27687 2485 27789
rect 12515 27687 12636 27789
rect 2364 27671 12636 27687
rect 13761 28894 13879 28928
rect 13761 28860 13801 28894
rect 13835 28860 13879 28894
rect 13761 28826 13879 28860
rect 13761 28792 13801 28826
rect 13835 28792 13879 28826
rect 13761 28758 13879 28792
rect 13761 28724 13801 28758
rect 13835 28724 13879 28758
rect 13761 28690 13879 28724
rect 13761 28656 13801 28690
rect 13835 28656 13879 28690
rect 13761 28622 13879 28656
rect 13761 28588 13801 28622
rect 13835 28588 13879 28622
rect 13761 28554 13879 28588
rect 13761 28520 13801 28554
rect 13835 28520 13879 28554
rect 13761 28486 13879 28520
rect 13761 28452 13801 28486
rect 13835 28452 13879 28486
rect 13761 28418 13879 28452
rect 13761 28384 13801 28418
rect 13835 28384 13879 28418
rect 13761 28350 13879 28384
rect 13761 28316 13801 28350
rect 13835 28316 13879 28350
rect 13761 28282 13879 28316
rect 13761 28248 13801 28282
rect 13835 28248 13879 28282
rect 13761 28214 13879 28248
rect 13761 28180 13801 28214
rect 13835 28180 13879 28214
rect 13761 28146 13879 28180
rect 13761 28112 13801 28146
rect 13835 28112 13879 28146
rect 13761 28078 13879 28112
rect 13761 28044 13801 28078
rect 13835 28044 13879 28078
rect 13761 28010 13879 28044
rect 13761 27976 13801 28010
rect 13835 27976 13879 28010
rect 13761 27942 13879 27976
rect 13761 27908 13801 27942
rect 13835 27908 13879 27942
rect 13761 27874 13879 27908
rect 13761 27840 13801 27874
rect 13835 27840 13879 27874
rect 13761 27806 13879 27840
rect 13761 27772 13801 27806
rect 13835 27772 13879 27806
rect 13761 27738 13879 27772
rect 13761 27704 13801 27738
rect 13835 27704 13879 27738
rect 13761 27670 13879 27704
rect 13761 27636 13801 27670
rect 13835 27636 13879 27670
rect 13761 27602 13879 27636
rect 13761 27568 13801 27602
rect 13835 27568 13879 27602
rect 13761 27534 13879 27568
rect 13761 27500 13801 27534
rect 13835 27500 13879 27534
rect 13761 27466 13879 27500
rect 13761 27432 13801 27466
rect 13835 27432 13879 27466
rect 13761 27398 13879 27432
rect 13761 27364 13801 27398
rect 13835 27364 13879 27398
rect 13761 27330 13879 27364
rect 13761 27296 13801 27330
rect 13835 27296 13879 27330
rect 13761 27262 13879 27296
rect 13761 27228 13801 27262
rect 13835 27228 13879 27262
rect 13761 27194 13879 27228
rect 13761 27160 13801 27194
rect 13835 27160 13879 27194
rect 13761 27126 13879 27160
rect 13761 27092 13801 27126
rect 13835 27092 13879 27126
rect 13761 27058 13879 27092
rect 1111 26995 1229 27029
rect 1111 26961 1153 26995
rect 1187 26961 1229 26995
rect 1111 26927 1229 26961
rect 1111 26893 1153 26927
rect 1187 26893 1229 26927
rect 1111 26859 1229 26893
rect 1111 26825 1153 26859
rect 1187 26825 1229 26859
rect 1111 26791 1229 26825
rect 1111 26757 1153 26791
rect 1187 26757 1229 26791
rect 1111 26723 1229 26757
rect 1111 26689 1153 26723
rect 1187 26689 1229 26723
rect 1111 26655 1229 26689
rect 1111 26621 1153 26655
rect 1187 26621 1229 26655
rect 1111 26587 1229 26621
rect 1111 26553 1153 26587
rect 1187 26553 1229 26587
rect 13761 27024 13801 27058
rect 13835 27024 13879 27058
rect 13761 26990 13879 27024
rect 13761 26956 13801 26990
rect 13835 26956 13879 26990
rect 13761 26922 13879 26956
rect 13761 26888 13801 26922
rect 13835 26888 13879 26922
rect 13761 26854 13879 26888
rect 13761 26820 13801 26854
rect 13835 26820 13879 26854
rect 13761 26786 13879 26820
rect 13761 26752 13801 26786
rect 13835 26752 13879 26786
rect 13761 26718 13879 26752
rect 13761 26684 13801 26718
rect 13835 26684 13879 26718
rect 13761 26650 13879 26684
rect 13761 26616 13801 26650
rect 13835 26616 13879 26650
rect 1111 26519 1229 26553
rect 1111 26485 1153 26519
rect 1187 26485 1229 26519
rect 1111 26451 1229 26485
rect 1111 26417 1153 26451
rect 1187 26417 1229 26451
rect 1111 26383 1229 26417
rect 1111 26349 1153 26383
rect 1187 26349 1229 26383
rect 1111 26315 1229 26349
rect 1111 26281 1153 26315
rect 1187 26281 1229 26315
rect 1111 26247 1229 26281
rect 1111 26213 1153 26247
rect 1187 26213 1229 26247
rect 1111 26179 1229 26213
rect 1111 26145 1153 26179
rect 1187 26145 1229 26179
rect 1111 26111 1229 26145
rect 1111 26077 1153 26111
rect 1187 26077 1229 26111
rect 1111 26043 1229 26077
rect 1111 26009 1153 26043
rect 1187 26009 1229 26043
rect 1111 25975 1229 26009
rect 1111 25941 1153 25975
rect 1187 25941 1229 25975
rect 1111 25907 1229 25941
rect 1111 25873 1153 25907
rect 1187 25873 1229 25907
rect 1111 25839 1229 25873
rect 1111 25805 1153 25839
rect 1187 25805 1229 25839
rect 1111 25771 1229 25805
rect 1111 25737 1153 25771
rect 1187 25737 1229 25771
rect 1111 25703 1229 25737
rect 1111 25669 1153 25703
rect 1187 25669 1229 25703
rect 1111 25635 1229 25669
rect 1111 25601 1153 25635
rect 1187 25601 1229 25635
rect 1111 25567 1229 25601
rect 1111 25533 1153 25567
rect 1187 25533 1229 25567
rect 1111 25499 1229 25533
rect 1111 25465 1153 25499
rect 1187 25465 1229 25499
rect 1111 25431 1229 25465
rect 1111 25397 1153 25431
rect 1187 25397 1229 25431
rect 1111 25363 1229 25397
rect 1111 25329 1153 25363
rect 1187 25329 1229 25363
rect 1111 25295 1229 25329
rect 1111 25261 1153 25295
rect 1187 25261 1229 25295
rect 1111 25227 1229 25261
rect 1111 25193 1153 25227
rect 1187 25193 1229 25227
rect 1111 25159 1229 25193
rect 1111 25125 1153 25159
rect 1187 25125 1229 25159
rect 1111 25091 1229 25125
rect 1111 25057 1153 25091
rect 1187 25057 1229 25091
rect 1111 25023 1229 25057
rect 1111 24989 1153 25023
rect 1187 24989 1229 25023
rect 1111 24955 1229 24989
rect 1111 24921 1153 24955
rect 1187 24921 1229 24955
rect 1111 24887 1229 24921
rect 1111 24853 1153 24887
rect 1187 24853 1229 24887
rect 1111 24819 1229 24853
rect 1748 26575 13228 26585
rect 1748 26201 2269 26575
rect 12707 26201 13228 26575
rect 1748 26191 13228 26201
rect 1748 26067 2142 26191
rect 1748 25353 1758 26067
rect 2132 25353 2142 26067
rect 12834 26067 13228 26191
rect 1748 25229 2142 25353
rect 12834 25353 12844 26067
rect 13218 25353 13228 26067
rect 12834 25229 13228 25353
rect 1748 25219 13228 25229
rect 1748 24845 2269 25219
rect 12707 24845 13228 25219
rect 1748 24835 13228 24845
rect 13761 26582 13879 26616
rect 13761 26548 13801 26582
rect 13835 26548 13879 26582
rect 13761 26514 13879 26548
rect 13761 26480 13801 26514
rect 13835 26480 13879 26514
rect 13761 26446 13879 26480
rect 13761 26412 13801 26446
rect 13835 26412 13879 26446
rect 13761 26378 13879 26412
rect 13761 26344 13801 26378
rect 13835 26344 13879 26378
rect 13761 26310 13879 26344
rect 13761 26276 13801 26310
rect 13835 26276 13879 26310
rect 13761 26242 13879 26276
rect 13761 26208 13801 26242
rect 13835 26208 13879 26242
rect 13761 26174 13879 26208
rect 13761 26140 13801 26174
rect 13835 26140 13879 26174
rect 13761 26106 13879 26140
rect 13761 26072 13801 26106
rect 13835 26072 13879 26106
rect 13761 26038 13879 26072
rect 13761 26004 13801 26038
rect 13835 26004 13879 26038
rect 13761 25970 13879 26004
rect 13761 25936 13801 25970
rect 13835 25936 13879 25970
rect 13761 25902 13879 25936
rect 13761 25868 13801 25902
rect 13835 25868 13879 25902
rect 13761 25834 13879 25868
rect 13761 25800 13801 25834
rect 13835 25800 13879 25834
rect 13761 25766 13879 25800
rect 13761 25732 13801 25766
rect 13835 25732 13879 25766
rect 13761 25698 13879 25732
rect 13761 25664 13801 25698
rect 13835 25664 13879 25698
rect 13761 25630 13879 25664
rect 13761 25596 13801 25630
rect 13835 25596 13879 25630
rect 13761 25562 13879 25596
rect 13761 25528 13801 25562
rect 13835 25528 13879 25562
rect 13761 25494 13879 25528
rect 13761 25460 13801 25494
rect 13835 25460 13879 25494
rect 13761 25426 13879 25460
rect 13761 25392 13801 25426
rect 13835 25392 13879 25426
rect 13761 25358 13879 25392
rect 13761 25324 13801 25358
rect 13835 25324 13879 25358
rect 13761 25290 13879 25324
rect 13761 25256 13801 25290
rect 13835 25256 13879 25290
rect 13761 25222 13879 25256
rect 13761 25188 13801 25222
rect 13835 25188 13879 25222
rect 13761 25154 13879 25188
rect 13761 25120 13801 25154
rect 13835 25120 13879 25154
rect 13761 25086 13879 25120
rect 13761 25052 13801 25086
rect 13835 25052 13879 25086
rect 13761 25018 13879 25052
rect 13761 24984 13801 25018
rect 13835 24984 13879 25018
rect 13761 24950 13879 24984
rect 13761 24916 13801 24950
rect 13835 24916 13879 24950
rect 13761 24882 13879 24916
rect 13761 24848 13801 24882
rect 13835 24848 13879 24882
rect 1111 24785 1153 24819
rect 1187 24785 1229 24819
rect 1111 24751 1229 24785
rect 1111 24717 1153 24751
rect 1187 24717 1229 24751
rect 1111 24683 1229 24717
rect 1111 24649 1153 24683
rect 1187 24649 1229 24683
rect 1111 24615 1229 24649
rect 1111 24581 1153 24615
rect 1187 24581 1229 24615
rect 1111 24547 1229 24581
rect 1111 24513 1153 24547
rect 1187 24513 1229 24547
rect 1111 24479 1229 24513
rect 1111 24445 1153 24479
rect 1187 24445 1229 24479
rect 1111 24411 1229 24445
rect 1111 24377 1153 24411
rect 1187 24377 1229 24411
rect 1111 24343 1229 24377
rect 1111 24309 1153 24343
rect 1187 24309 1229 24343
rect 1111 24275 1229 24309
rect 1111 24241 1153 24275
rect 1187 24241 1229 24275
rect 1111 24207 1229 24241
rect 1111 24173 1153 24207
rect 1187 24173 1229 24207
rect 1111 24139 1229 24173
rect 1111 24105 1153 24139
rect 1187 24105 1229 24139
rect 1111 24071 1229 24105
rect 1111 24037 1153 24071
rect 1187 24037 1229 24071
rect 1111 24003 1229 24037
rect 1111 23969 1153 24003
rect 1187 23969 1229 24003
rect 1111 23935 1229 23969
rect 1111 23901 1153 23935
rect 1187 23901 1229 23935
rect 1111 23867 1229 23901
rect 1111 23833 1153 23867
rect 1187 23833 1229 23867
rect 1111 23799 1229 23833
rect 1111 23765 1153 23799
rect 1187 23765 1229 23799
rect 1111 23731 1229 23765
rect 1111 23697 1153 23731
rect 1187 23697 1229 23731
rect 1111 23663 1229 23697
rect 1111 23629 1153 23663
rect 1187 23629 1229 23663
rect 1111 23595 1229 23629
rect 1111 23561 1153 23595
rect 1187 23561 1229 23595
rect 1111 23527 1229 23561
rect 1111 23493 1153 23527
rect 1187 23493 1229 23527
rect 1111 23459 1229 23493
rect 1111 23425 1153 23459
rect 1187 23425 1229 23459
rect 1111 23391 1229 23425
rect 1111 23357 1153 23391
rect 1187 23357 1229 23391
rect 1111 23323 1229 23357
rect 1111 23289 1153 23323
rect 1187 23289 1229 23323
rect 1111 23255 1229 23289
rect 1111 23221 1153 23255
rect 1187 23221 1229 23255
rect 1111 23187 1229 23221
rect 1111 23153 1153 23187
rect 1187 23153 1229 23187
rect 1111 23119 1229 23153
rect 1111 23085 1153 23119
rect 1187 23085 1229 23119
rect 1111 23051 1229 23085
rect 1111 23017 1153 23051
rect 1187 23017 1229 23051
rect 1111 22983 1229 23017
rect 1111 22949 1153 22983
rect 1187 22949 1229 22983
rect 1111 22915 1229 22949
rect 1111 22881 1153 22915
rect 1187 22881 1229 22915
rect 1111 22847 1229 22881
rect 1111 22813 1153 22847
rect 1187 22813 1229 22847
rect 1111 22779 1229 22813
rect 1111 22745 1153 22779
rect 1187 22745 1229 22779
rect 1111 22711 1229 22745
rect 1111 22677 1153 22711
rect 1187 22677 1229 22711
rect 1111 22643 1229 22677
rect 1111 22609 1153 22643
rect 1187 22609 1229 22643
rect 1111 22575 1229 22609
rect 1111 22541 1153 22575
rect 1187 22541 1229 22575
rect 1111 22507 1229 22541
rect 1111 22473 1153 22507
rect 1187 22473 1229 22507
rect 1111 22439 1229 22473
rect 1111 22405 1153 22439
rect 1187 22405 1229 22439
rect 1111 22371 1229 22405
rect 1111 22337 1153 22371
rect 1187 22337 1229 22371
rect 1111 22303 1229 22337
rect 1111 22269 1153 22303
rect 1187 22269 1229 22303
rect 1111 22235 1229 22269
rect 1111 22201 1153 22235
rect 1187 22201 1229 22235
rect 1111 22167 1229 22201
rect 1111 22133 1153 22167
rect 1187 22133 1229 22167
rect 1111 22099 1229 22133
rect 1111 22065 1153 22099
rect 1187 22065 1229 22099
rect 1111 22031 1229 22065
rect 1111 21997 1153 22031
rect 1187 21997 1229 22031
rect 1111 21963 1229 21997
rect 1111 21929 1153 21963
rect 1187 21929 1229 21963
rect 1111 21895 1229 21929
rect 1111 21861 1153 21895
rect 1187 21861 1229 21895
rect 1111 21827 1229 21861
rect 1111 21793 1153 21827
rect 1187 21793 1229 21827
rect 1111 21759 1229 21793
rect 1111 21725 1153 21759
rect 1187 21725 1229 21759
rect 1111 21691 1229 21725
rect 1111 21657 1153 21691
rect 1187 21657 1229 21691
rect 1111 21623 1229 21657
rect 1111 21589 1153 21623
rect 1187 21589 1229 21623
rect 1111 21555 1229 21589
rect 1111 21521 1153 21555
rect 1187 21521 1229 21555
rect 1111 21487 1229 21521
rect 1111 21453 1153 21487
rect 1187 21453 1229 21487
rect 1111 21419 1229 21453
rect 1111 21385 1153 21419
rect 1187 21385 1229 21419
rect 1111 21351 1229 21385
rect 1111 21317 1153 21351
rect 1187 21317 1229 21351
rect 1111 21283 1229 21317
rect 1111 21249 1153 21283
rect 1187 21249 1229 21283
rect 1111 21215 1229 21249
rect 1111 21181 1153 21215
rect 1187 21181 1229 21215
rect 1111 21147 1229 21181
rect 1111 21113 1153 21147
rect 1187 21113 1229 21147
rect 1111 21079 1229 21113
rect 1111 21045 1153 21079
rect 1187 21045 1229 21079
rect 1111 21011 1229 21045
rect 1111 20977 1153 21011
rect 1187 20977 1229 21011
rect 1111 20943 1229 20977
rect 1111 20909 1153 20943
rect 1187 20909 1229 20943
rect 1111 20875 1229 20909
rect 1111 20841 1153 20875
rect 1187 20841 1229 20875
rect 1111 20807 1229 20841
rect 1111 20773 1153 20807
rect 1187 20773 1229 20807
rect 1111 20739 1229 20773
rect 1111 20705 1153 20739
rect 1187 20705 1229 20739
rect 1111 20671 1229 20705
rect 1111 20637 1153 20671
rect 1187 20637 1229 20671
rect 1111 20603 1229 20637
rect 1111 20569 1153 20603
rect 1187 20569 1229 20603
rect 1111 20535 1229 20569
rect 1111 20501 1153 20535
rect 1187 20501 1229 20535
rect 1111 20467 1229 20501
rect 1111 20433 1153 20467
rect 1187 20433 1229 20467
rect 1111 20399 1229 20433
rect 1111 20365 1153 20399
rect 1187 20365 1229 20399
rect 1111 20331 1229 20365
rect 1111 20297 1153 20331
rect 1187 20297 1229 20331
rect 1111 20263 1229 20297
rect 1111 20229 1153 20263
rect 1187 20229 1229 20263
rect 1111 20195 1229 20229
rect 1111 20161 1153 20195
rect 1187 20161 1229 20195
rect 1111 20127 1229 20161
rect 1111 20093 1153 20127
rect 1187 20093 1229 20127
rect 1111 20059 1229 20093
rect 1111 20025 1153 20059
rect 1187 20025 1229 20059
rect 1111 19991 1229 20025
rect 1111 19957 1153 19991
rect 1187 19957 1229 19991
rect 1111 19923 1229 19957
rect 1111 19889 1153 19923
rect 1187 19889 1229 19923
rect 1111 19855 1229 19889
rect 1111 19821 1153 19855
rect 1187 19821 1229 19855
rect 1111 19787 1229 19821
rect 1111 19753 1153 19787
rect 1187 19753 1229 19787
rect 1111 19719 1229 19753
rect 1111 19685 1153 19719
rect 1187 19685 1229 19719
rect 1111 19651 1229 19685
rect 1111 19617 1153 19651
rect 1187 19617 1229 19651
rect 1111 19583 1229 19617
rect 1111 19549 1153 19583
rect 1187 19549 1229 19583
rect 1111 19515 1229 19549
rect 1111 19481 1153 19515
rect 1187 19481 1229 19515
rect 1111 19447 1229 19481
rect 1111 19413 1153 19447
rect 1187 19413 1229 19447
rect 1111 19379 1229 19413
rect 1111 19345 1153 19379
rect 1187 19345 1229 19379
rect 1111 19311 1229 19345
rect 1111 19277 1153 19311
rect 1187 19277 1229 19311
rect 1111 19243 1229 19277
rect 1111 19209 1153 19243
rect 1187 19209 1229 19243
rect 1111 19175 1229 19209
rect 1111 19141 1153 19175
rect 1187 19141 1229 19175
rect 1111 19107 1229 19141
rect 1111 19073 1153 19107
rect 1187 19073 1229 19107
rect 1111 19039 1229 19073
rect 1111 19005 1153 19039
rect 1187 19005 1229 19039
rect 1111 18971 1229 19005
rect 1111 18937 1153 18971
rect 1187 18937 1229 18971
rect 1111 18903 1229 18937
rect 1111 18869 1153 18903
rect 1187 18869 1229 18903
rect 1111 18835 1229 18869
rect 1111 18801 1153 18835
rect 1187 18801 1229 18835
rect 1111 18767 1229 18801
rect 1111 18733 1153 18767
rect 1187 18733 1229 18767
rect 1111 18699 1229 18733
rect 1111 18665 1153 18699
rect 1187 18665 1229 18699
rect 1111 18631 1229 18665
rect 1111 18597 1153 18631
rect 1187 18597 1229 18631
rect 1111 18563 1229 18597
rect 1111 18529 1153 18563
rect 1187 18529 1229 18563
rect 1111 18495 1229 18529
rect 1111 18461 1153 18495
rect 1187 18461 1229 18495
rect 1111 18427 1229 18461
rect 1111 18393 1153 18427
rect 1187 18393 1229 18427
rect 1111 18359 1229 18393
rect 1111 18325 1153 18359
rect 1187 18325 1229 18359
rect 1111 18291 1229 18325
rect 1111 18257 1153 18291
rect 1187 18257 1229 18291
rect 1111 18223 1229 18257
rect 1111 18189 1153 18223
rect 1187 18189 1229 18223
rect 1111 18155 1229 18189
rect 1111 18121 1153 18155
rect 1187 18121 1229 18155
rect 1111 18087 1229 18121
rect 1111 18053 1153 18087
rect 1187 18053 1229 18087
rect 1111 18019 1229 18053
rect 1111 17985 1153 18019
rect 1187 17985 1229 18019
rect 1111 17951 1229 17985
rect 1111 17917 1153 17951
rect 1187 17917 1229 17951
rect 1111 17883 1229 17917
rect 1111 17849 1153 17883
rect 1187 17849 1229 17883
rect 1111 17815 1229 17849
rect 1111 17781 1153 17815
rect 1187 17781 1229 17815
rect 1111 17747 1229 17781
rect 1111 17713 1153 17747
rect 1187 17713 1229 17747
rect 1111 17679 1229 17713
rect 1111 17645 1153 17679
rect 1187 17645 1229 17679
rect 1111 17611 1229 17645
rect 1111 17577 1153 17611
rect 1187 17577 1229 17611
rect 1111 17543 1229 17577
rect 1111 17509 1153 17543
rect 1187 17509 1229 17543
rect 1111 17475 1229 17509
rect 1111 17441 1153 17475
rect 1187 17441 1229 17475
rect 1111 17407 1229 17441
rect 1111 17373 1153 17407
rect 1187 17373 1229 17407
rect 1111 17339 1229 17373
rect 1111 17305 1153 17339
rect 1187 17305 1229 17339
rect 1111 17271 1229 17305
rect 1111 17237 1153 17271
rect 1187 17237 1229 17271
rect 1111 17203 1229 17237
rect 1111 17169 1153 17203
rect 1187 17169 1229 17203
rect 1111 17135 1229 17169
rect 1111 17101 1153 17135
rect 1187 17101 1229 17135
rect 1111 17067 1229 17101
rect 1111 17033 1153 17067
rect 1187 17033 1229 17067
rect 1111 16999 1229 17033
rect 1111 16965 1153 16999
rect 1187 16965 1229 16999
rect 1111 16931 1229 16965
rect 1111 16897 1153 16931
rect 1187 16897 1229 16931
rect 1111 16863 1229 16897
rect 1111 16829 1153 16863
rect 1187 16829 1229 16863
rect 1111 16795 1229 16829
rect 1111 16761 1153 16795
rect 1187 16761 1229 16795
rect 1111 16727 1229 16761
rect 1111 16693 1153 16727
rect 1187 16693 1229 16727
rect 1111 16659 1229 16693
rect 1111 16625 1153 16659
rect 1187 16625 1229 16659
rect 1111 16591 1229 16625
rect 1111 16557 1153 16591
rect 1187 16557 1229 16591
rect 1111 16523 1229 16557
rect 1111 16489 1153 16523
rect 1187 16489 1229 16523
rect 1111 16455 1229 16489
rect 1111 16421 1153 16455
rect 1187 16421 1229 16455
rect 1111 16387 1229 16421
rect 1111 16353 1153 16387
rect 1187 16353 1229 16387
rect 1111 16319 1229 16353
rect 1111 16285 1153 16319
rect 1187 16285 1229 16319
rect 1111 16251 1229 16285
rect 1111 16217 1153 16251
rect 1187 16217 1229 16251
rect 1111 16183 1229 16217
rect 1111 16149 1153 16183
rect 1187 16149 1229 16183
rect 1111 16115 1229 16149
rect 1111 16081 1153 16115
rect 1187 16081 1229 16115
rect 1111 16047 1229 16081
rect 1111 16013 1153 16047
rect 1187 16013 1229 16047
rect 1111 15979 1229 16013
rect 1111 15945 1153 15979
rect 1187 15945 1229 15979
rect 1111 15911 1229 15945
rect 1111 15877 1153 15911
rect 1187 15877 1229 15911
rect 1111 15843 1229 15877
rect 1111 15809 1153 15843
rect 1187 15809 1229 15843
rect 1111 15775 1229 15809
rect 1111 15741 1153 15775
rect 1187 15741 1229 15775
rect 1111 15707 1229 15741
rect 1111 15673 1153 15707
rect 1187 15673 1229 15707
rect 1111 15639 1229 15673
rect 1111 15605 1153 15639
rect 1187 15605 1229 15639
rect 1111 15571 1229 15605
rect 1111 15537 1153 15571
rect 1187 15537 1229 15571
rect 1111 15503 1229 15537
rect 1111 15469 1153 15503
rect 1187 15469 1229 15503
rect 1111 15435 1229 15469
rect 1111 15401 1153 15435
rect 1187 15401 1229 15435
rect 1111 15332 1229 15401
rect 13761 24814 13879 24848
rect 13761 24780 13801 24814
rect 13835 24780 13879 24814
rect 13761 24746 13879 24780
rect 13761 24712 13801 24746
rect 13835 24712 13879 24746
rect 13761 24678 13879 24712
rect 13761 24644 13801 24678
rect 13835 24644 13879 24678
rect 13761 24610 13879 24644
rect 13761 24576 13801 24610
rect 13835 24576 13879 24610
rect 13761 24542 13879 24576
rect 13761 24508 13801 24542
rect 13835 24508 13879 24542
rect 13761 24474 13879 24508
rect 13761 24440 13801 24474
rect 13835 24440 13879 24474
rect 13761 24406 13879 24440
rect 13761 24372 13801 24406
rect 13835 24372 13879 24406
rect 13761 24338 13879 24372
rect 13761 24304 13801 24338
rect 13835 24304 13879 24338
rect 13761 24270 13879 24304
rect 13761 24236 13801 24270
rect 13835 24236 13879 24270
rect 13761 24202 13879 24236
rect 13761 24168 13801 24202
rect 13835 24168 13879 24202
rect 13761 24134 13879 24168
rect 13761 24100 13801 24134
rect 13835 24100 13879 24134
rect 13761 24066 13879 24100
rect 13761 24032 13801 24066
rect 13835 24032 13879 24066
rect 13761 23998 13879 24032
rect 13761 23964 13801 23998
rect 13835 23964 13879 23998
rect 13761 23930 13879 23964
rect 13761 23896 13801 23930
rect 13835 23896 13879 23930
rect 13761 23862 13879 23896
rect 13761 23828 13801 23862
rect 13835 23828 13879 23862
rect 13761 23794 13879 23828
rect 13761 23760 13801 23794
rect 13835 23760 13879 23794
rect 13761 23726 13879 23760
rect 13761 23692 13801 23726
rect 13835 23692 13879 23726
rect 13761 23658 13879 23692
rect 13761 23624 13801 23658
rect 13835 23624 13879 23658
rect 13761 23590 13879 23624
rect 13761 23556 13801 23590
rect 13835 23556 13879 23590
rect 13761 23522 13879 23556
rect 13761 23488 13801 23522
rect 13835 23488 13879 23522
rect 13761 23454 13879 23488
rect 13761 23420 13801 23454
rect 13835 23420 13879 23454
rect 13761 23386 13879 23420
rect 13761 23352 13801 23386
rect 13835 23352 13879 23386
rect 13761 23318 13879 23352
rect 13761 23284 13801 23318
rect 13835 23284 13879 23318
rect 13761 23250 13879 23284
rect 13761 23216 13801 23250
rect 13835 23216 13879 23250
rect 13761 23182 13879 23216
rect 13761 23148 13801 23182
rect 13835 23148 13879 23182
rect 13761 23114 13879 23148
rect 13761 23080 13801 23114
rect 13835 23080 13879 23114
rect 13761 23046 13879 23080
rect 13761 23012 13801 23046
rect 13835 23012 13879 23046
rect 13761 22978 13879 23012
rect 13761 22944 13801 22978
rect 13835 22944 13879 22978
rect 13761 22910 13879 22944
rect 13761 22876 13801 22910
rect 13835 22876 13879 22910
rect 13761 22842 13879 22876
rect 13761 22808 13801 22842
rect 13835 22808 13879 22842
rect 13761 22774 13879 22808
rect 13761 22740 13801 22774
rect 13835 22740 13879 22774
rect 13761 22706 13879 22740
rect 13761 22672 13801 22706
rect 13835 22672 13879 22706
rect 13761 22638 13879 22672
rect 13761 22604 13801 22638
rect 13835 22604 13879 22638
rect 13761 22570 13879 22604
rect 13761 22536 13801 22570
rect 13835 22536 13879 22570
rect 13761 22502 13879 22536
rect 13761 22468 13801 22502
rect 13835 22468 13879 22502
rect 13761 22434 13879 22468
rect 13761 22400 13801 22434
rect 13835 22400 13879 22434
rect 13761 22366 13879 22400
rect 13761 22332 13801 22366
rect 13835 22332 13879 22366
rect 13761 22298 13879 22332
rect 13761 22264 13801 22298
rect 13835 22264 13879 22298
rect 13761 22230 13879 22264
rect 13761 22196 13801 22230
rect 13835 22196 13879 22230
rect 13761 22162 13879 22196
rect 13761 22128 13801 22162
rect 13835 22128 13879 22162
rect 13761 22094 13879 22128
rect 13761 22060 13801 22094
rect 13835 22060 13879 22094
rect 13761 22026 13879 22060
rect 13761 21992 13801 22026
rect 13835 21992 13879 22026
rect 13761 21958 13879 21992
rect 13761 21924 13801 21958
rect 13835 21924 13879 21958
rect 13761 21890 13879 21924
rect 13761 21856 13801 21890
rect 13835 21856 13879 21890
rect 13761 21822 13879 21856
rect 13761 21788 13801 21822
rect 13835 21788 13879 21822
rect 13761 21754 13879 21788
rect 13761 21720 13801 21754
rect 13835 21720 13879 21754
rect 13761 21686 13879 21720
rect 13761 21652 13801 21686
rect 13835 21652 13879 21686
rect 13761 21618 13879 21652
rect 13761 21584 13801 21618
rect 13835 21584 13879 21618
rect 13761 21550 13879 21584
rect 13761 21516 13801 21550
rect 13835 21516 13879 21550
rect 13761 21482 13879 21516
rect 13761 21448 13801 21482
rect 13835 21448 13879 21482
rect 13761 21414 13879 21448
rect 13761 21380 13801 21414
rect 13835 21380 13879 21414
rect 13761 21346 13879 21380
rect 13761 21312 13801 21346
rect 13835 21312 13879 21346
rect 13761 21278 13879 21312
rect 13761 21244 13801 21278
rect 13835 21244 13879 21278
rect 13761 21210 13879 21244
rect 13761 21176 13801 21210
rect 13835 21176 13879 21210
rect 13761 21142 13879 21176
rect 13761 21108 13801 21142
rect 13835 21108 13879 21142
rect 13761 21074 13879 21108
rect 13761 21040 13801 21074
rect 13835 21040 13879 21074
rect 13761 21006 13879 21040
rect 13761 20972 13801 21006
rect 13835 20972 13879 21006
rect 13761 20938 13879 20972
rect 13761 20904 13801 20938
rect 13835 20904 13879 20938
rect 13761 20870 13879 20904
rect 13761 20836 13801 20870
rect 13835 20836 13879 20870
rect 13761 20802 13879 20836
rect 13761 20768 13801 20802
rect 13835 20768 13879 20802
rect 13761 20734 13879 20768
rect 13761 20700 13801 20734
rect 13835 20700 13879 20734
rect 13761 20666 13879 20700
rect 13761 20632 13801 20666
rect 13835 20632 13879 20666
rect 13761 20598 13879 20632
rect 13761 20564 13801 20598
rect 13835 20564 13879 20598
rect 13761 20530 13879 20564
rect 13761 20496 13801 20530
rect 13835 20496 13879 20530
rect 13761 20462 13879 20496
rect 13761 20428 13801 20462
rect 13835 20428 13879 20462
rect 13761 20394 13879 20428
rect 13761 20360 13801 20394
rect 13835 20360 13879 20394
rect 13761 20326 13879 20360
rect 13761 20292 13801 20326
rect 13835 20292 13879 20326
rect 13761 20258 13879 20292
rect 13761 20224 13801 20258
rect 13835 20224 13879 20258
rect 13761 20190 13879 20224
rect 13761 20156 13801 20190
rect 13835 20156 13879 20190
rect 13761 20122 13879 20156
rect 13761 20088 13801 20122
rect 13835 20088 13879 20122
rect 13761 20054 13879 20088
rect 13761 20020 13801 20054
rect 13835 20020 13879 20054
rect 13761 19986 13879 20020
rect 13761 19952 13801 19986
rect 13835 19952 13879 19986
rect 13761 19918 13879 19952
rect 13761 19884 13801 19918
rect 13835 19884 13879 19918
rect 13761 19850 13879 19884
rect 13761 19816 13801 19850
rect 13835 19816 13879 19850
rect 13761 19782 13879 19816
rect 13761 19748 13801 19782
rect 13835 19748 13879 19782
rect 13761 19714 13879 19748
rect 13761 19680 13801 19714
rect 13835 19680 13879 19714
rect 13761 19646 13879 19680
rect 13761 19612 13801 19646
rect 13835 19612 13879 19646
rect 13761 19578 13879 19612
rect 13761 19544 13801 19578
rect 13835 19544 13879 19578
rect 13761 19510 13879 19544
rect 13761 19476 13801 19510
rect 13835 19476 13879 19510
rect 13761 19442 13879 19476
rect 13761 19408 13801 19442
rect 13835 19408 13879 19442
rect 13761 19374 13879 19408
rect 13761 19340 13801 19374
rect 13835 19340 13879 19374
rect 13761 19306 13879 19340
rect 13761 19272 13801 19306
rect 13835 19272 13879 19306
rect 13761 19238 13879 19272
rect 13761 19204 13801 19238
rect 13835 19204 13879 19238
rect 13761 19170 13879 19204
rect 13761 19136 13801 19170
rect 13835 19136 13879 19170
rect 13761 19102 13879 19136
rect 13761 19068 13801 19102
rect 13835 19068 13879 19102
rect 13761 19034 13879 19068
rect 13761 19000 13801 19034
rect 13835 19000 13879 19034
rect 13761 18966 13879 19000
rect 13761 18932 13801 18966
rect 13835 18932 13879 18966
rect 13761 18898 13879 18932
rect 13761 18864 13801 18898
rect 13835 18864 13879 18898
rect 13761 18830 13879 18864
rect 13761 18796 13801 18830
rect 13835 18796 13879 18830
rect 13761 18762 13879 18796
rect 13761 18728 13801 18762
rect 13835 18728 13879 18762
rect 13761 18694 13879 18728
rect 13761 18660 13801 18694
rect 13835 18660 13879 18694
rect 13761 18626 13879 18660
rect 13761 18592 13801 18626
rect 13835 18592 13879 18626
rect 13761 18558 13879 18592
rect 13761 18524 13801 18558
rect 13835 18524 13879 18558
rect 13761 18490 13879 18524
rect 13761 18456 13801 18490
rect 13835 18456 13879 18490
rect 13761 18422 13879 18456
rect 13761 18388 13801 18422
rect 13835 18388 13879 18422
rect 13761 18354 13879 18388
rect 13761 18320 13801 18354
rect 13835 18320 13879 18354
rect 13761 18286 13879 18320
rect 13761 18252 13801 18286
rect 13835 18252 13879 18286
rect 13761 18218 13879 18252
rect 13761 18184 13801 18218
rect 13835 18184 13879 18218
rect 13761 18150 13879 18184
rect 13761 18116 13801 18150
rect 13835 18116 13879 18150
rect 13761 18082 13879 18116
rect 13761 18048 13801 18082
rect 13835 18048 13879 18082
rect 13761 18014 13879 18048
rect 13761 17980 13801 18014
rect 13835 17980 13879 18014
rect 13761 17946 13879 17980
rect 13761 17912 13801 17946
rect 13835 17912 13879 17946
rect 13761 17878 13879 17912
rect 13761 17844 13801 17878
rect 13835 17844 13879 17878
rect 13761 17810 13879 17844
rect 13761 17776 13801 17810
rect 13835 17776 13879 17810
rect 13761 17742 13879 17776
rect 13761 17708 13801 17742
rect 13835 17708 13879 17742
rect 13761 17674 13879 17708
rect 13761 17640 13801 17674
rect 13835 17640 13879 17674
rect 13761 17606 13879 17640
rect 13761 17572 13801 17606
rect 13835 17572 13879 17606
rect 13761 17538 13879 17572
rect 13761 17504 13801 17538
rect 13835 17504 13879 17538
rect 13761 17470 13879 17504
rect 13761 17436 13801 17470
rect 13835 17436 13879 17470
rect 13761 17402 13879 17436
rect 13761 17368 13801 17402
rect 13835 17368 13879 17402
rect 13761 17334 13879 17368
rect 13761 17300 13801 17334
rect 13835 17300 13879 17334
rect 13761 17266 13879 17300
rect 13761 17232 13801 17266
rect 13835 17232 13879 17266
rect 13761 17198 13879 17232
rect 13761 17164 13801 17198
rect 13835 17164 13879 17198
rect 13761 17130 13879 17164
rect 13761 17096 13801 17130
rect 13835 17096 13879 17130
rect 13761 17062 13879 17096
rect 13761 17028 13801 17062
rect 13835 17028 13879 17062
rect 13761 16994 13879 17028
rect 13761 16960 13801 16994
rect 13835 16960 13879 16994
rect 13761 16926 13879 16960
rect 13761 16892 13801 16926
rect 13835 16892 13879 16926
rect 13761 16858 13879 16892
rect 13761 16824 13801 16858
rect 13835 16824 13879 16858
rect 13761 16790 13879 16824
rect 13761 16756 13801 16790
rect 13835 16756 13879 16790
rect 13761 16722 13879 16756
rect 13761 16688 13801 16722
rect 13835 16688 13879 16722
rect 13761 16654 13879 16688
rect 13761 16620 13801 16654
rect 13835 16620 13879 16654
rect 13761 16586 13879 16620
rect 13761 16552 13801 16586
rect 13835 16552 13879 16586
rect 13761 16518 13879 16552
rect 13761 16484 13801 16518
rect 13835 16484 13879 16518
rect 13761 16450 13879 16484
rect 13761 16416 13801 16450
rect 13835 16416 13879 16450
rect 13761 16382 13879 16416
rect 13761 16348 13801 16382
rect 13835 16348 13879 16382
rect 13761 16314 13879 16348
rect 13761 16280 13801 16314
rect 13835 16280 13879 16314
rect 13761 16246 13879 16280
rect 13761 16212 13801 16246
rect 13835 16212 13879 16246
rect 13761 16178 13879 16212
rect 13761 16144 13801 16178
rect 13835 16144 13879 16178
rect 13761 16110 13879 16144
rect 13761 16076 13801 16110
rect 13835 16076 13879 16110
rect 13761 16042 13879 16076
rect 13761 16008 13801 16042
rect 13835 16008 13879 16042
rect 13761 15974 13879 16008
rect 13761 15940 13801 15974
rect 13835 15940 13879 15974
rect 13761 15906 13879 15940
rect 13761 15872 13801 15906
rect 13835 15872 13879 15906
rect 13761 15838 13879 15872
rect 13761 15804 13801 15838
rect 13835 15804 13879 15838
rect 13761 15770 13879 15804
rect 13761 15736 13801 15770
rect 13835 15736 13879 15770
rect 13761 15702 13879 15736
rect 13761 15668 13801 15702
rect 13835 15668 13879 15702
rect 13761 15634 13879 15668
rect 13761 15600 13801 15634
rect 13835 15600 13879 15634
rect 13761 15566 13879 15600
rect 13761 15532 13801 15566
rect 13835 15532 13879 15566
rect 13761 15498 13879 15532
rect 13761 15464 13801 15498
rect 13835 15464 13879 15498
rect 13761 15430 13879 15464
rect 13761 15396 13801 15430
rect 13835 15396 13879 15430
rect 13761 15332 13879 15396
rect 1111 15291 13879 15332
rect 1111 15257 1294 15291
rect 1328 15257 1362 15291
rect 1396 15257 1430 15291
rect 1464 15257 1498 15291
rect 1532 15257 1566 15291
rect 1600 15257 1634 15291
rect 1668 15257 1702 15291
rect 1736 15257 1770 15291
rect 1804 15257 1838 15291
rect 1872 15257 1906 15291
rect 1940 15257 1974 15291
rect 2008 15257 2042 15291
rect 2076 15257 2110 15291
rect 2144 15257 2178 15291
rect 2212 15257 2246 15291
rect 2280 15257 2314 15291
rect 2348 15257 2382 15291
rect 2416 15257 2450 15291
rect 2484 15257 2518 15291
rect 2552 15257 2586 15291
rect 2620 15257 2654 15291
rect 2688 15257 2722 15291
rect 2756 15257 2790 15291
rect 2824 15257 2858 15291
rect 2892 15257 2926 15291
rect 2960 15257 2994 15291
rect 3028 15257 3062 15291
rect 3096 15257 3130 15291
rect 3164 15257 3198 15291
rect 3232 15257 3266 15291
rect 3300 15257 3334 15291
rect 3368 15257 3402 15291
rect 3436 15257 3470 15291
rect 3504 15257 3538 15291
rect 3572 15257 3606 15291
rect 3640 15257 3674 15291
rect 3708 15257 3742 15291
rect 3776 15257 3810 15291
rect 3844 15257 3878 15291
rect 3912 15257 3946 15291
rect 3980 15257 4014 15291
rect 4048 15257 4082 15291
rect 4116 15257 4150 15291
rect 4184 15257 4218 15291
rect 4252 15257 4286 15291
rect 4320 15257 4354 15291
rect 4388 15257 4422 15291
rect 4456 15257 4490 15291
rect 4524 15257 4558 15291
rect 4592 15257 4626 15291
rect 4660 15257 4694 15291
rect 4728 15257 4762 15291
rect 4796 15257 4830 15291
rect 4864 15257 4898 15291
rect 4932 15257 4966 15291
rect 5000 15257 5034 15291
rect 5068 15257 5102 15291
rect 5136 15257 5170 15291
rect 5204 15257 5238 15291
rect 5272 15257 5306 15291
rect 5340 15257 5374 15291
rect 5408 15257 5442 15291
rect 5476 15257 5510 15291
rect 5544 15257 5578 15291
rect 5612 15257 5646 15291
rect 5680 15257 5714 15291
rect 5748 15257 5782 15291
rect 5816 15257 5850 15291
rect 5884 15257 5918 15291
rect 5952 15257 5986 15291
rect 6020 15257 6054 15291
rect 6088 15257 6122 15291
rect 6156 15257 6190 15291
rect 6224 15257 6258 15291
rect 6292 15257 6326 15291
rect 6360 15257 6394 15291
rect 6428 15257 6462 15291
rect 6496 15257 6530 15291
rect 6564 15257 6598 15291
rect 6632 15257 6666 15291
rect 6700 15257 6734 15291
rect 6768 15257 6802 15291
rect 6836 15257 6870 15291
rect 6904 15257 6938 15291
rect 6972 15257 7006 15291
rect 7040 15257 7074 15291
rect 7108 15257 7142 15291
rect 7176 15257 7210 15291
rect 7244 15257 7278 15291
rect 7312 15257 7346 15291
rect 7380 15257 7414 15291
rect 7448 15257 7482 15291
rect 7516 15257 7550 15291
rect 7584 15257 7618 15291
rect 7652 15257 7686 15291
rect 7720 15257 7754 15291
rect 7788 15257 7822 15291
rect 7856 15257 7890 15291
rect 7924 15257 7958 15291
rect 7992 15257 8026 15291
rect 8060 15257 8094 15291
rect 8128 15257 8162 15291
rect 8196 15257 8230 15291
rect 8264 15257 8298 15291
rect 8332 15257 8366 15291
rect 8400 15257 8434 15291
rect 8468 15257 8502 15291
rect 8536 15257 8570 15291
rect 8604 15257 8638 15291
rect 8672 15257 8706 15291
rect 8740 15257 8774 15291
rect 8808 15257 8842 15291
rect 8876 15257 8910 15291
rect 8944 15257 8978 15291
rect 9012 15257 9046 15291
rect 9080 15257 9114 15291
rect 9148 15257 9182 15291
rect 9216 15257 9250 15291
rect 9284 15257 9318 15291
rect 9352 15257 9386 15291
rect 9420 15257 9454 15291
rect 9488 15257 9522 15291
rect 9556 15257 9590 15291
rect 9624 15257 9658 15291
rect 9692 15257 9726 15291
rect 9760 15257 9794 15291
rect 9828 15257 9862 15291
rect 9896 15257 9930 15291
rect 9964 15257 9998 15291
rect 10032 15257 10066 15291
rect 10100 15257 10134 15291
rect 10168 15257 10202 15291
rect 10236 15257 10270 15291
rect 10304 15257 10338 15291
rect 10372 15257 10406 15291
rect 10440 15257 10474 15291
rect 10508 15257 10542 15291
rect 10576 15257 10610 15291
rect 10644 15257 10678 15291
rect 10712 15257 10746 15291
rect 10780 15257 10814 15291
rect 10848 15257 10882 15291
rect 10916 15257 10950 15291
rect 10984 15257 11018 15291
rect 11052 15257 11086 15291
rect 11120 15257 11154 15291
rect 11188 15257 11222 15291
rect 11256 15257 11290 15291
rect 11324 15257 11358 15291
rect 11392 15257 11426 15291
rect 11460 15257 11494 15291
rect 11528 15257 11562 15291
rect 11596 15257 11630 15291
rect 11664 15257 11698 15291
rect 11732 15257 11766 15291
rect 11800 15257 11834 15291
rect 11868 15257 11902 15291
rect 11936 15257 11970 15291
rect 12004 15257 12038 15291
rect 12072 15257 12106 15291
rect 12140 15257 12174 15291
rect 12208 15257 12242 15291
rect 12276 15257 12310 15291
rect 12344 15257 12378 15291
rect 12412 15257 12446 15291
rect 12480 15257 12514 15291
rect 12548 15257 12582 15291
rect 12616 15257 12650 15291
rect 12684 15257 12718 15291
rect 12752 15257 12786 15291
rect 12820 15257 12854 15291
rect 12888 15257 12922 15291
rect 12956 15257 12990 15291
rect 13024 15257 13058 15291
rect 13092 15257 13126 15291
rect 13160 15257 13194 15291
rect 13228 15257 13262 15291
rect 13296 15257 13330 15291
rect 13364 15257 13398 15291
rect 13432 15257 13466 15291
rect 13500 15257 13534 15291
rect 13568 15257 13602 15291
rect 13636 15257 13670 15291
rect 13704 15257 13879 15291
rect 1111 15214 13879 15257
rect 14531 36239 14716 36273
rect 14531 36205 14599 36239
rect 14633 36205 14716 36239
rect 14531 36171 14716 36205
rect 14531 36137 14599 36171
rect 14633 36137 14716 36171
rect 14531 36103 14716 36137
rect 14531 36069 14599 36103
rect 14633 36069 14716 36103
rect 14531 36035 14716 36069
rect 14531 36001 14599 36035
rect 14633 36001 14716 36035
rect 14531 35967 14716 36001
rect 14531 35933 14599 35967
rect 14633 35933 14716 35967
rect 14531 35899 14716 35933
rect 14531 35865 14599 35899
rect 14633 35865 14716 35899
rect 14531 35831 14716 35865
rect 14531 35797 14599 35831
rect 14633 35797 14716 35831
rect 14531 35763 14716 35797
rect 14531 35729 14599 35763
rect 14633 35729 14716 35763
rect 14531 35695 14716 35729
rect 14531 35661 14599 35695
rect 14633 35661 14716 35695
rect 14531 35627 14716 35661
rect 14531 35593 14599 35627
rect 14633 35593 14716 35627
rect 14531 35559 14716 35593
rect 14531 35525 14599 35559
rect 14633 35525 14716 35559
rect 14531 35491 14716 35525
rect 14531 35457 14599 35491
rect 14633 35457 14716 35491
rect 14531 35423 14716 35457
rect 14531 35389 14599 35423
rect 14633 35389 14716 35423
rect 14531 35355 14716 35389
rect 14531 35321 14599 35355
rect 14633 35321 14716 35355
rect 14531 35287 14716 35321
rect 14531 35253 14599 35287
rect 14633 35253 14716 35287
rect 14531 35219 14716 35253
rect 14531 35185 14599 35219
rect 14633 35185 14716 35219
rect 14531 35151 14716 35185
rect 14531 35117 14599 35151
rect 14633 35117 14716 35151
rect 14531 35083 14716 35117
rect 14531 35049 14599 35083
rect 14633 35049 14716 35083
rect 14531 35015 14716 35049
rect 14531 34981 14599 35015
rect 14633 34981 14716 35015
rect 14531 34947 14716 34981
rect 14531 34913 14599 34947
rect 14633 34913 14716 34947
rect 14531 34879 14716 34913
rect 14531 34845 14599 34879
rect 14633 34845 14716 34879
rect 14531 34811 14716 34845
rect 14531 34777 14599 34811
rect 14633 34777 14716 34811
rect 14531 34743 14716 34777
rect 14531 34709 14599 34743
rect 14633 34709 14716 34743
rect 14531 34675 14716 34709
rect 14531 34641 14599 34675
rect 14633 34641 14716 34675
rect 14531 34607 14716 34641
rect 14531 34573 14599 34607
rect 14633 34573 14716 34607
rect 14531 34539 14716 34573
rect 14531 34505 14599 34539
rect 14633 34505 14716 34539
rect 14531 34471 14716 34505
rect 14531 34437 14599 34471
rect 14633 34437 14716 34471
rect 14531 34403 14716 34437
rect 14531 34369 14599 34403
rect 14633 34369 14716 34403
rect 14531 34335 14716 34369
rect 14531 34301 14599 34335
rect 14633 34301 14716 34335
rect 14531 34267 14716 34301
rect 14531 34233 14599 34267
rect 14633 34233 14716 34267
rect 14531 34199 14716 34233
rect 14531 34165 14599 34199
rect 14633 34165 14716 34199
rect 14531 34131 14716 34165
rect 14531 34097 14599 34131
rect 14633 34097 14716 34131
rect 14531 34063 14716 34097
rect 14531 34029 14599 34063
rect 14633 34029 14716 34063
rect 14531 33995 14716 34029
rect 14531 33961 14599 33995
rect 14633 33961 14716 33995
rect 14531 33927 14716 33961
rect 14531 33893 14599 33927
rect 14633 33893 14716 33927
rect 14531 33859 14716 33893
rect 14531 33825 14599 33859
rect 14633 33825 14716 33859
rect 14531 33791 14716 33825
rect 14531 33757 14599 33791
rect 14633 33757 14716 33791
rect 14531 33723 14716 33757
rect 14531 33689 14599 33723
rect 14633 33689 14716 33723
rect 14531 33655 14716 33689
rect 14531 33621 14599 33655
rect 14633 33621 14716 33655
rect 14531 33587 14716 33621
rect 14531 33553 14599 33587
rect 14633 33553 14716 33587
rect 14531 33519 14716 33553
rect 14531 33485 14599 33519
rect 14633 33485 14716 33519
rect 14531 33451 14716 33485
rect 14531 33417 14599 33451
rect 14633 33417 14716 33451
rect 14531 33383 14716 33417
rect 14531 33349 14599 33383
rect 14633 33349 14716 33383
rect 14531 33315 14716 33349
rect 14531 33281 14599 33315
rect 14633 33281 14716 33315
rect 14531 33247 14716 33281
rect 14531 33213 14599 33247
rect 14633 33213 14716 33247
rect 14531 33179 14716 33213
rect 14531 33145 14599 33179
rect 14633 33145 14716 33179
rect 14531 33111 14716 33145
rect 14531 33077 14599 33111
rect 14633 33077 14716 33111
rect 14531 33043 14716 33077
rect 14531 33009 14599 33043
rect 14633 33009 14716 33043
rect 14531 32975 14716 33009
rect 14531 32941 14599 32975
rect 14633 32941 14716 32975
rect 14531 32907 14716 32941
rect 14531 32873 14599 32907
rect 14633 32873 14716 32907
rect 14531 32839 14716 32873
rect 14531 32805 14599 32839
rect 14633 32805 14716 32839
rect 14531 32771 14716 32805
rect 14531 32737 14599 32771
rect 14633 32737 14716 32771
rect 14531 32703 14716 32737
rect 14531 32669 14599 32703
rect 14633 32669 14716 32703
rect 14531 32635 14716 32669
rect 14531 32601 14599 32635
rect 14633 32601 14716 32635
rect 14531 32567 14716 32601
rect 14531 32533 14599 32567
rect 14633 32533 14716 32567
rect 14531 32499 14716 32533
rect 14531 32465 14599 32499
rect 14633 32465 14716 32499
rect 14531 32431 14716 32465
rect 14531 32397 14599 32431
rect 14633 32397 14716 32431
rect 14531 32363 14716 32397
rect 14531 32329 14599 32363
rect 14633 32329 14716 32363
rect 14531 32295 14716 32329
rect 14531 32261 14599 32295
rect 14633 32261 14716 32295
rect 14531 32227 14716 32261
rect 14531 32193 14599 32227
rect 14633 32193 14716 32227
rect 14531 32159 14716 32193
rect 14531 32125 14599 32159
rect 14633 32125 14716 32159
rect 14531 32091 14716 32125
rect 14531 32057 14599 32091
rect 14633 32057 14716 32091
rect 14531 32023 14716 32057
rect 14531 31989 14599 32023
rect 14633 31989 14716 32023
rect 14531 31955 14716 31989
rect 14531 31921 14599 31955
rect 14633 31921 14716 31955
rect 14531 31887 14716 31921
rect 14531 31853 14599 31887
rect 14633 31853 14716 31887
rect 14531 31819 14716 31853
rect 14531 31785 14599 31819
rect 14633 31785 14716 31819
rect 14531 31751 14716 31785
rect 14531 31717 14599 31751
rect 14633 31717 14716 31751
rect 14531 31683 14716 31717
rect 14531 31649 14599 31683
rect 14633 31649 14716 31683
rect 14531 31615 14716 31649
rect 14531 31581 14599 31615
rect 14633 31581 14716 31615
rect 14531 31547 14716 31581
rect 14531 31513 14599 31547
rect 14633 31513 14716 31547
rect 14531 31479 14716 31513
rect 14531 31445 14599 31479
rect 14633 31445 14716 31479
rect 14531 31411 14716 31445
rect 14531 31377 14599 31411
rect 14633 31377 14716 31411
rect 14531 31343 14716 31377
rect 14531 31309 14599 31343
rect 14633 31309 14716 31343
rect 14531 31275 14716 31309
rect 14531 31241 14599 31275
rect 14633 31241 14716 31275
rect 14531 31207 14716 31241
rect 14531 31173 14599 31207
rect 14633 31173 14716 31207
rect 14531 31139 14716 31173
rect 14531 31105 14599 31139
rect 14633 31105 14716 31139
rect 14531 31071 14716 31105
rect 14531 31037 14599 31071
rect 14633 31037 14716 31071
rect 14531 31003 14716 31037
rect 14531 30969 14599 31003
rect 14633 30969 14716 31003
rect 14531 30935 14716 30969
rect 14531 30901 14599 30935
rect 14633 30901 14716 30935
rect 14531 30867 14716 30901
rect 14531 30833 14599 30867
rect 14633 30833 14716 30867
rect 14531 30799 14716 30833
rect 14531 30765 14599 30799
rect 14633 30765 14716 30799
rect 14531 30731 14716 30765
rect 14531 30697 14599 30731
rect 14633 30697 14716 30731
rect 14531 30663 14716 30697
rect 14531 30629 14599 30663
rect 14633 30629 14716 30663
rect 14531 30595 14716 30629
rect 14531 30561 14599 30595
rect 14633 30561 14716 30595
rect 14531 30527 14716 30561
rect 14531 30493 14599 30527
rect 14633 30493 14716 30527
rect 14531 30459 14716 30493
rect 14531 30425 14599 30459
rect 14633 30425 14716 30459
rect 14531 30391 14716 30425
rect 14531 30357 14599 30391
rect 14633 30357 14716 30391
rect 14531 30323 14716 30357
rect 14531 30289 14599 30323
rect 14633 30289 14716 30323
rect 14531 30255 14716 30289
rect 14531 30221 14599 30255
rect 14633 30221 14716 30255
rect 14531 30187 14716 30221
rect 14531 30153 14599 30187
rect 14633 30153 14716 30187
rect 14531 30119 14716 30153
rect 14531 30085 14599 30119
rect 14633 30085 14716 30119
rect 14531 30051 14716 30085
rect 14531 30017 14599 30051
rect 14633 30017 14716 30051
rect 14531 29983 14716 30017
rect 14531 29949 14599 29983
rect 14633 29949 14716 29983
rect 14531 29915 14716 29949
rect 14531 29881 14599 29915
rect 14633 29881 14716 29915
rect 14531 29847 14716 29881
rect 14531 29813 14599 29847
rect 14633 29813 14716 29847
rect 14531 29779 14716 29813
rect 14531 29745 14599 29779
rect 14633 29745 14716 29779
rect 14531 29711 14716 29745
rect 14531 29677 14599 29711
rect 14633 29677 14716 29711
rect 14531 29643 14716 29677
rect 14531 29609 14599 29643
rect 14633 29609 14716 29643
rect 14531 29575 14716 29609
rect 14531 29541 14599 29575
rect 14633 29541 14716 29575
rect 14531 29507 14716 29541
rect 14531 29473 14599 29507
rect 14633 29473 14716 29507
rect 14531 29439 14716 29473
rect 14531 29405 14599 29439
rect 14633 29405 14716 29439
rect 14531 29371 14716 29405
rect 14531 29337 14599 29371
rect 14633 29337 14716 29371
rect 14531 29303 14716 29337
rect 14531 29269 14599 29303
rect 14633 29269 14716 29303
rect 14531 29235 14716 29269
rect 14531 29201 14599 29235
rect 14633 29201 14716 29235
rect 14531 29167 14716 29201
rect 14531 29133 14599 29167
rect 14633 29133 14716 29167
rect 14531 29099 14716 29133
rect 14531 29065 14599 29099
rect 14633 29065 14716 29099
rect 14531 29031 14716 29065
rect 14531 28997 14599 29031
rect 14633 28997 14716 29031
rect 14531 28963 14716 28997
rect 14531 28929 14599 28963
rect 14633 28929 14716 28963
rect 14531 28895 14716 28929
rect 14531 28861 14599 28895
rect 14633 28861 14716 28895
rect 14531 28827 14716 28861
rect 14531 28793 14599 28827
rect 14633 28793 14716 28827
rect 14531 28759 14716 28793
rect 14531 28725 14599 28759
rect 14633 28725 14716 28759
rect 14531 28691 14716 28725
rect 14531 28657 14599 28691
rect 14633 28657 14716 28691
rect 14531 28623 14716 28657
rect 14531 28589 14599 28623
rect 14633 28589 14716 28623
rect 14531 28555 14716 28589
rect 14531 28521 14599 28555
rect 14633 28521 14716 28555
rect 14531 28487 14716 28521
rect 14531 28453 14599 28487
rect 14633 28453 14716 28487
rect 14531 28419 14716 28453
rect 14531 28385 14599 28419
rect 14633 28385 14716 28419
rect 14531 28351 14716 28385
rect 14531 28317 14599 28351
rect 14633 28317 14716 28351
rect 14531 28283 14716 28317
rect 14531 28249 14599 28283
rect 14633 28249 14716 28283
rect 14531 28215 14716 28249
rect 14531 28181 14599 28215
rect 14633 28181 14716 28215
rect 14531 28147 14716 28181
rect 14531 28113 14599 28147
rect 14633 28113 14716 28147
rect 14531 28079 14716 28113
rect 14531 28045 14599 28079
rect 14633 28045 14716 28079
rect 14531 28011 14716 28045
rect 14531 27977 14599 28011
rect 14633 27977 14716 28011
rect 14531 27943 14716 27977
rect 14531 27909 14599 27943
rect 14633 27909 14716 27943
rect 14531 27875 14716 27909
rect 14531 27841 14599 27875
rect 14633 27841 14716 27875
rect 14531 27807 14716 27841
rect 14531 27773 14599 27807
rect 14633 27773 14716 27807
rect 14531 27739 14716 27773
rect 14531 27705 14599 27739
rect 14633 27705 14716 27739
rect 14531 27671 14716 27705
rect 14531 27637 14599 27671
rect 14633 27637 14716 27671
rect 14531 27603 14716 27637
rect 14531 27569 14599 27603
rect 14633 27569 14716 27603
rect 14531 27535 14716 27569
rect 14531 27501 14599 27535
rect 14633 27501 14716 27535
rect 14531 27467 14716 27501
rect 14531 27433 14599 27467
rect 14633 27433 14716 27467
rect 14531 27399 14716 27433
rect 14531 27365 14599 27399
rect 14633 27365 14716 27399
rect 14531 27331 14716 27365
rect 14531 27297 14599 27331
rect 14633 27297 14716 27331
rect 14531 27263 14716 27297
rect 14531 27229 14599 27263
rect 14633 27229 14716 27263
rect 14531 27195 14716 27229
rect 14531 27161 14599 27195
rect 14633 27161 14716 27195
rect 14531 27127 14716 27161
rect 14531 27093 14599 27127
rect 14633 27093 14716 27127
rect 14531 27059 14716 27093
rect 14531 27025 14599 27059
rect 14633 27025 14716 27059
rect 14531 26991 14716 27025
rect 14531 26957 14599 26991
rect 14633 26957 14716 26991
rect 14531 26923 14716 26957
rect 14531 26889 14599 26923
rect 14633 26889 14716 26923
rect 14531 26855 14716 26889
rect 14531 26821 14599 26855
rect 14633 26821 14716 26855
rect 14531 26787 14716 26821
rect 14531 26753 14599 26787
rect 14633 26753 14716 26787
rect 14531 26719 14716 26753
rect 14531 26685 14599 26719
rect 14633 26685 14716 26719
rect 14531 26651 14716 26685
rect 14531 26617 14599 26651
rect 14633 26617 14716 26651
rect 14531 26583 14716 26617
rect 14531 26549 14599 26583
rect 14633 26549 14716 26583
rect 14531 26515 14716 26549
rect 14531 26481 14599 26515
rect 14633 26481 14716 26515
rect 14531 26447 14716 26481
rect 14531 26413 14599 26447
rect 14633 26413 14716 26447
rect 14531 26379 14716 26413
rect 14531 26345 14599 26379
rect 14633 26345 14716 26379
rect 14531 26311 14716 26345
rect 14531 26277 14599 26311
rect 14633 26277 14716 26311
rect 14531 26243 14716 26277
rect 14531 26209 14599 26243
rect 14633 26209 14716 26243
rect 14531 26175 14716 26209
rect 14531 26141 14599 26175
rect 14633 26141 14716 26175
rect 14531 26107 14716 26141
rect 14531 26073 14599 26107
rect 14633 26073 14716 26107
rect 14531 26039 14716 26073
rect 14531 26005 14599 26039
rect 14633 26005 14716 26039
rect 14531 25971 14716 26005
rect 14531 25937 14599 25971
rect 14633 25937 14716 25971
rect 14531 25903 14716 25937
rect 14531 25869 14599 25903
rect 14633 25869 14716 25903
rect 14531 25835 14716 25869
rect 14531 25801 14599 25835
rect 14633 25801 14716 25835
rect 14531 25767 14716 25801
rect 14531 25733 14599 25767
rect 14633 25733 14716 25767
rect 14531 25699 14716 25733
rect 14531 25665 14599 25699
rect 14633 25665 14716 25699
rect 14531 25631 14716 25665
rect 14531 25597 14599 25631
rect 14633 25597 14716 25631
rect 14531 25563 14716 25597
rect 14531 25529 14599 25563
rect 14633 25529 14716 25563
rect 14531 25495 14716 25529
rect 14531 25461 14599 25495
rect 14633 25461 14716 25495
rect 14531 25427 14716 25461
rect 14531 25393 14599 25427
rect 14633 25393 14716 25427
rect 14531 25359 14716 25393
rect 14531 25325 14599 25359
rect 14633 25325 14716 25359
rect 14531 25291 14716 25325
rect 14531 25257 14599 25291
rect 14633 25257 14716 25291
rect 14531 25223 14716 25257
rect 14531 25189 14599 25223
rect 14633 25189 14716 25223
rect 14531 25155 14716 25189
rect 14531 25121 14599 25155
rect 14633 25121 14716 25155
rect 14531 25087 14716 25121
rect 14531 25053 14599 25087
rect 14633 25053 14716 25087
rect 14531 25019 14716 25053
rect 14531 24985 14599 25019
rect 14633 24985 14716 25019
rect 14531 24951 14716 24985
rect 14531 24917 14599 24951
rect 14633 24917 14716 24951
rect 14531 24883 14716 24917
rect 14531 24849 14599 24883
rect 14633 24849 14716 24883
rect 14531 24815 14716 24849
rect 14531 24781 14599 24815
rect 14633 24781 14716 24815
rect 14531 24747 14716 24781
rect 14531 24713 14599 24747
rect 14633 24713 14716 24747
rect 14531 24679 14716 24713
rect 14531 24645 14599 24679
rect 14633 24645 14716 24679
rect 14531 24611 14716 24645
rect 14531 24577 14599 24611
rect 14633 24577 14716 24611
rect 14531 24543 14716 24577
rect 14531 24509 14599 24543
rect 14633 24509 14716 24543
rect 14531 24475 14716 24509
rect 14531 24441 14599 24475
rect 14633 24441 14716 24475
rect 14531 24407 14716 24441
rect 14531 24373 14599 24407
rect 14633 24373 14716 24407
rect 14531 24339 14716 24373
rect 14531 24305 14599 24339
rect 14633 24305 14716 24339
rect 14531 24271 14716 24305
rect 14531 24237 14599 24271
rect 14633 24237 14716 24271
rect 14531 24203 14716 24237
rect 14531 24169 14599 24203
rect 14633 24169 14716 24203
rect 14531 24135 14716 24169
rect 14531 24101 14599 24135
rect 14633 24101 14716 24135
rect 14531 24067 14716 24101
rect 14531 24033 14599 24067
rect 14633 24033 14716 24067
rect 14531 23999 14716 24033
rect 14531 23965 14599 23999
rect 14633 23965 14716 23999
rect 14531 23931 14716 23965
rect 14531 23897 14599 23931
rect 14633 23897 14716 23931
rect 14531 23863 14716 23897
rect 14531 23829 14599 23863
rect 14633 23829 14716 23863
rect 14531 23795 14716 23829
rect 14531 23761 14599 23795
rect 14633 23761 14716 23795
rect 14531 23727 14716 23761
rect 14531 23693 14599 23727
rect 14633 23693 14716 23727
rect 14531 23659 14716 23693
rect 14531 23625 14599 23659
rect 14633 23625 14716 23659
rect 14531 23591 14716 23625
rect 14531 23557 14599 23591
rect 14633 23557 14716 23591
rect 14531 23523 14716 23557
rect 14531 23489 14599 23523
rect 14633 23489 14716 23523
rect 14531 23455 14716 23489
rect 14531 23421 14599 23455
rect 14633 23421 14716 23455
rect 14531 23387 14716 23421
rect 14531 23353 14599 23387
rect 14633 23353 14716 23387
rect 14531 23319 14716 23353
rect 14531 23285 14599 23319
rect 14633 23285 14716 23319
rect 14531 23251 14716 23285
rect 14531 23217 14599 23251
rect 14633 23217 14716 23251
rect 14531 23183 14716 23217
rect 14531 23149 14599 23183
rect 14633 23149 14716 23183
rect 14531 23115 14716 23149
rect 14531 23081 14599 23115
rect 14633 23081 14716 23115
rect 14531 23047 14716 23081
rect 14531 23013 14599 23047
rect 14633 23013 14716 23047
rect 14531 22979 14716 23013
rect 14531 22945 14599 22979
rect 14633 22945 14716 22979
rect 14531 22911 14716 22945
rect 14531 22877 14599 22911
rect 14633 22877 14716 22911
rect 14531 22843 14716 22877
rect 14531 22809 14599 22843
rect 14633 22809 14716 22843
rect 14531 22775 14716 22809
rect 14531 22741 14599 22775
rect 14633 22741 14716 22775
rect 14531 22707 14716 22741
rect 14531 22673 14599 22707
rect 14633 22673 14716 22707
rect 14531 22639 14716 22673
rect 14531 22605 14599 22639
rect 14633 22605 14716 22639
rect 14531 22571 14716 22605
rect 14531 22537 14599 22571
rect 14633 22537 14716 22571
rect 14531 22503 14716 22537
rect 14531 22469 14599 22503
rect 14633 22469 14716 22503
rect 14531 22435 14716 22469
rect 14531 22401 14599 22435
rect 14633 22401 14716 22435
rect 14531 22367 14716 22401
rect 14531 22333 14599 22367
rect 14633 22333 14716 22367
rect 14531 22299 14716 22333
rect 14531 22265 14599 22299
rect 14633 22265 14716 22299
rect 14531 22231 14716 22265
rect 14531 22197 14599 22231
rect 14633 22197 14716 22231
rect 14531 22163 14716 22197
rect 14531 22129 14599 22163
rect 14633 22129 14716 22163
rect 14531 22095 14716 22129
rect 14531 22061 14599 22095
rect 14633 22061 14716 22095
rect 14531 22027 14716 22061
rect 14531 21993 14599 22027
rect 14633 21993 14716 22027
rect 14531 21959 14716 21993
rect 14531 21925 14599 21959
rect 14633 21925 14716 21959
rect 14531 21891 14716 21925
rect 14531 21857 14599 21891
rect 14633 21857 14716 21891
rect 14531 21823 14716 21857
rect 14531 21789 14599 21823
rect 14633 21789 14716 21823
rect 14531 21755 14716 21789
rect 14531 21721 14599 21755
rect 14633 21721 14716 21755
rect 14531 21687 14716 21721
rect 14531 21653 14599 21687
rect 14633 21653 14716 21687
rect 14531 21619 14716 21653
rect 14531 21585 14599 21619
rect 14633 21585 14716 21619
rect 14531 21551 14716 21585
rect 14531 21517 14599 21551
rect 14633 21517 14716 21551
rect 14531 21483 14716 21517
rect 14531 21449 14599 21483
rect 14633 21449 14716 21483
rect 14531 21415 14716 21449
rect 14531 21381 14599 21415
rect 14633 21381 14716 21415
rect 14531 21347 14716 21381
rect 14531 21313 14599 21347
rect 14633 21313 14716 21347
rect 14531 21279 14716 21313
rect 14531 21245 14599 21279
rect 14633 21245 14716 21279
rect 14531 21211 14716 21245
rect 14531 21177 14599 21211
rect 14633 21177 14716 21211
rect 14531 21143 14716 21177
rect 14531 21109 14599 21143
rect 14633 21109 14716 21143
rect 14531 21075 14716 21109
rect 14531 21041 14599 21075
rect 14633 21041 14716 21075
rect 14531 21007 14716 21041
rect 14531 20973 14599 21007
rect 14633 20973 14716 21007
rect 14531 20939 14716 20973
rect 14531 20905 14599 20939
rect 14633 20905 14716 20939
rect 14531 20871 14716 20905
rect 14531 20837 14599 20871
rect 14633 20837 14716 20871
rect 14531 20803 14716 20837
rect 14531 20769 14599 20803
rect 14633 20769 14716 20803
rect 14531 20735 14716 20769
rect 14531 20701 14599 20735
rect 14633 20701 14716 20735
rect 14531 20667 14716 20701
rect 14531 20633 14599 20667
rect 14633 20633 14716 20667
rect 14531 20599 14716 20633
rect 14531 20565 14599 20599
rect 14633 20565 14716 20599
rect 14531 20531 14716 20565
rect 14531 20497 14599 20531
rect 14633 20497 14716 20531
rect 14531 20463 14716 20497
rect 14531 20429 14599 20463
rect 14633 20429 14716 20463
rect 14531 20395 14716 20429
rect 14531 20361 14599 20395
rect 14633 20361 14716 20395
rect 14531 20327 14716 20361
rect 14531 20293 14599 20327
rect 14633 20293 14716 20327
rect 14531 20259 14716 20293
rect 14531 20225 14599 20259
rect 14633 20225 14716 20259
rect 14531 20191 14716 20225
rect 14531 20157 14599 20191
rect 14633 20157 14716 20191
rect 14531 20123 14716 20157
rect 14531 20089 14599 20123
rect 14633 20089 14716 20123
rect 14531 20055 14716 20089
rect 14531 20021 14599 20055
rect 14633 20021 14716 20055
rect 14531 19987 14716 20021
rect 14531 19953 14599 19987
rect 14633 19953 14716 19987
rect 14531 19919 14716 19953
rect 14531 19885 14599 19919
rect 14633 19885 14716 19919
rect 14531 19851 14716 19885
rect 14531 19817 14599 19851
rect 14633 19817 14716 19851
rect 14531 19783 14716 19817
rect 14531 19749 14599 19783
rect 14633 19749 14716 19783
rect 14531 19715 14716 19749
rect 14531 19681 14599 19715
rect 14633 19681 14716 19715
rect 14531 19647 14716 19681
rect 14531 19613 14599 19647
rect 14633 19613 14716 19647
rect 14531 19579 14716 19613
rect 14531 19545 14599 19579
rect 14633 19545 14716 19579
rect 14531 19511 14716 19545
rect 14531 19477 14599 19511
rect 14633 19477 14716 19511
rect 14531 19443 14716 19477
rect 14531 19409 14599 19443
rect 14633 19409 14716 19443
rect 14531 19375 14716 19409
rect 14531 19341 14599 19375
rect 14633 19341 14716 19375
rect 14531 19307 14716 19341
rect 14531 19273 14599 19307
rect 14633 19273 14716 19307
rect 14531 19239 14716 19273
rect 14531 19205 14599 19239
rect 14633 19205 14716 19239
rect 14531 19171 14716 19205
rect 14531 19137 14599 19171
rect 14633 19137 14716 19171
rect 14531 19103 14716 19137
rect 14531 19069 14599 19103
rect 14633 19069 14716 19103
rect 14531 19035 14716 19069
rect 14531 19001 14599 19035
rect 14633 19001 14716 19035
rect 14531 18967 14716 19001
rect 14531 18933 14599 18967
rect 14633 18933 14716 18967
rect 14531 18899 14716 18933
rect 14531 18865 14599 18899
rect 14633 18865 14716 18899
rect 14531 18831 14716 18865
rect 14531 18797 14599 18831
rect 14633 18797 14716 18831
rect 14531 18763 14716 18797
rect 14531 18729 14599 18763
rect 14633 18729 14716 18763
rect 14531 18695 14716 18729
rect 14531 18661 14599 18695
rect 14633 18661 14716 18695
rect 14531 18627 14716 18661
rect 14531 18593 14599 18627
rect 14633 18593 14716 18627
rect 14531 18559 14716 18593
rect 14531 18525 14599 18559
rect 14633 18525 14716 18559
rect 14531 18491 14716 18525
rect 14531 18457 14599 18491
rect 14633 18457 14716 18491
rect 14531 18423 14716 18457
rect 14531 18389 14599 18423
rect 14633 18389 14716 18423
rect 14531 18355 14716 18389
rect 14531 18321 14599 18355
rect 14633 18321 14716 18355
rect 14531 18287 14716 18321
rect 14531 18253 14599 18287
rect 14633 18253 14716 18287
rect 14531 18219 14716 18253
rect 14531 18185 14599 18219
rect 14633 18185 14716 18219
rect 14531 18151 14716 18185
rect 14531 18117 14599 18151
rect 14633 18117 14716 18151
rect 14531 18083 14716 18117
rect 14531 18049 14599 18083
rect 14633 18049 14716 18083
rect 14531 18015 14716 18049
rect 14531 17981 14599 18015
rect 14633 17981 14716 18015
rect 14531 17947 14716 17981
rect 14531 17913 14599 17947
rect 14633 17913 14716 17947
rect 14531 17879 14716 17913
rect 14531 17845 14599 17879
rect 14633 17845 14716 17879
rect 14531 17811 14716 17845
rect 14531 17777 14599 17811
rect 14633 17777 14716 17811
rect 14531 17743 14716 17777
rect 14531 17709 14599 17743
rect 14633 17709 14716 17743
rect 14531 17675 14716 17709
rect 14531 17641 14599 17675
rect 14633 17641 14716 17675
rect 14531 17607 14716 17641
rect 14531 17573 14599 17607
rect 14633 17573 14716 17607
rect 14531 17539 14716 17573
rect 14531 17505 14599 17539
rect 14633 17505 14716 17539
rect 14531 17471 14716 17505
rect 14531 17437 14599 17471
rect 14633 17437 14716 17471
rect 14531 17403 14716 17437
rect 14531 17369 14599 17403
rect 14633 17369 14716 17403
rect 14531 17335 14716 17369
rect 14531 17301 14599 17335
rect 14633 17301 14716 17335
rect 14531 17267 14716 17301
rect 14531 17233 14599 17267
rect 14633 17233 14716 17267
rect 14531 17199 14716 17233
rect 14531 17165 14599 17199
rect 14633 17165 14716 17199
rect 14531 17131 14716 17165
rect 14531 17097 14599 17131
rect 14633 17097 14716 17131
rect 14531 17063 14716 17097
rect 14531 17029 14599 17063
rect 14633 17029 14716 17063
rect 14531 16995 14716 17029
rect 14531 16961 14599 16995
rect 14633 16961 14716 16995
rect 14531 16927 14716 16961
rect 14531 16893 14599 16927
rect 14633 16893 14716 16927
rect 14531 16859 14716 16893
rect 14531 16825 14599 16859
rect 14633 16825 14716 16859
rect 14531 16791 14716 16825
rect 14531 16757 14599 16791
rect 14633 16757 14716 16791
rect 14531 16723 14716 16757
rect 14531 16689 14599 16723
rect 14633 16689 14716 16723
rect 14531 16655 14716 16689
rect 14531 16621 14599 16655
rect 14633 16621 14716 16655
rect 14531 16587 14716 16621
rect 14531 16553 14599 16587
rect 14633 16553 14716 16587
rect 14531 16519 14716 16553
rect 14531 16485 14599 16519
rect 14633 16485 14716 16519
rect 14531 16451 14716 16485
rect 14531 16417 14599 16451
rect 14633 16417 14716 16451
rect 14531 16383 14716 16417
rect 14531 16349 14599 16383
rect 14633 16349 14716 16383
rect 14531 16315 14716 16349
rect 14531 16281 14599 16315
rect 14633 16281 14716 16315
rect 14531 16247 14716 16281
rect 14531 16213 14599 16247
rect 14633 16213 14716 16247
rect 14531 16179 14716 16213
rect 14531 16145 14599 16179
rect 14633 16145 14716 16179
rect 14531 16111 14716 16145
rect 14531 16077 14599 16111
rect 14633 16077 14716 16111
rect 14531 16043 14716 16077
rect 14531 16009 14599 16043
rect 14633 16009 14716 16043
rect 14531 15975 14716 16009
rect 14531 15941 14599 15975
rect 14633 15941 14716 15975
rect 14531 15907 14716 15941
rect 14531 15873 14599 15907
rect 14633 15873 14716 15907
rect 14531 15839 14716 15873
rect 14531 15805 14599 15839
rect 14633 15805 14716 15839
rect 14531 15771 14716 15805
rect 14531 15737 14599 15771
rect 14633 15737 14716 15771
rect 14531 15703 14716 15737
rect 14531 15669 14599 15703
rect 14633 15669 14716 15703
rect 14531 15635 14716 15669
rect 14531 15601 14599 15635
rect 14633 15601 14716 15635
rect 14531 15567 14716 15601
rect 14531 15533 14599 15567
rect 14633 15533 14716 15567
rect 14531 15499 14716 15533
rect 14531 15465 14599 15499
rect 14633 15465 14716 15499
rect 14531 15431 14716 15465
rect 14531 15397 14599 15431
rect 14633 15397 14716 15431
rect 14531 15363 14716 15397
rect 14531 15329 14599 15363
rect 14633 15329 14716 15363
rect 14531 15295 14716 15329
rect 14531 15261 14599 15295
rect 14633 15261 14716 15295
rect 14531 15227 14716 15261
rect 14531 15193 14599 15227
rect 14633 15193 14716 15227
rect 14531 15159 14716 15193
rect 14531 15125 14599 15159
rect 14633 15125 14716 15159
rect 14531 15091 14716 15125
rect 14531 15057 14599 15091
rect 14633 15057 14716 15091
rect 14531 15023 14716 15057
rect 14531 14989 14599 15023
rect 14633 14989 14716 15023
rect 14531 14955 14716 14989
rect 14531 14921 14599 14955
rect 14633 14921 14716 14955
rect 14531 14887 14716 14921
rect 14531 14853 14599 14887
rect 14633 14853 14716 14887
rect 14531 14819 14716 14853
rect 14531 14785 14599 14819
rect 14633 14785 14716 14819
rect 14531 14751 14716 14785
rect 14531 14717 14599 14751
rect 14633 14717 14716 14751
rect 237 14643 304 14677
rect 338 14643 422 14677
rect 237 14609 422 14643
rect 237 14575 304 14609
rect 338 14575 422 14609
rect 237 14541 422 14575
rect 14531 14683 14716 14717
rect 14531 14649 14599 14683
rect 14633 14649 14716 14683
rect 14531 14615 14716 14649
rect 14531 14581 14599 14615
rect 14633 14581 14716 14615
rect 14531 14541 14716 14581
rect 237 14464 14716 14541
rect 237 14430 468 14464
rect 502 14430 536 14464
rect 570 14430 604 14464
rect 638 14430 672 14464
rect 706 14430 740 14464
rect 774 14430 808 14464
rect 842 14430 876 14464
rect 910 14430 944 14464
rect 978 14430 1012 14464
rect 1046 14430 1080 14464
rect 1114 14430 1148 14464
rect 1182 14430 1216 14464
rect 1250 14430 1284 14464
rect 1318 14430 1352 14464
rect 1386 14430 1420 14464
rect 1454 14430 1488 14464
rect 1522 14430 1556 14464
rect 1590 14430 1624 14464
rect 1658 14430 1692 14464
rect 1726 14430 1760 14464
rect 1794 14430 1828 14464
rect 1862 14430 1896 14464
rect 1930 14430 1964 14464
rect 1998 14430 2032 14464
rect 2066 14430 2100 14464
rect 2134 14430 2168 14464
rect 2202 14430 2236 14464
rect 2270 14430 2304 14464
rect 2338 14430 2372 14464
rect 2406 14430 2440 14464
rect 2474 14430 2508 14464
rect 2542 14430 2576 14464
rect 2610 14430 2644 14464
rect 2678 14430 2712 14464
rect 2746 14430 2780 14464
rect 2814 14430 2848 14464
rect 2882 14430 2916 14464
rect 2950 14430 2984 14464
rect 3018 14430 3052 14464
rect 3086 14430 3120 14464
rect 3154 14430 3188 14464
rect 3222 14430 3256 14464
rect 3290 14430 3324 14464
rect 3358 14430 3392 14464
rect 3426 14430 3460 14464
rect 3494 14430 3528 14464
rect 3562 14430 3596 14464
rect 3630 14430 3664 14464
rect 3698 14430 3732 14464
rect 3766 14430 3800 14464
rect 3834 14430 3868 14464
rect 3902 14430 3936 14464
rect 3970 14430 4004 14464
rect 4038 14430 4072 14464
rect 4106 14430 4140 14464
rect 4174 14430 4208 14464
rect 4242 14430 4276 14464
rect 4310 14430 4344 14464
rect 4378 14430 4412 14464
rect 4446 14430 4480 14464
rect 4514 14430 4548 14464
rect 4582 14430 4616 14464
rect 4650 14430 4684 14464
rect 4718 14430 4752 14464
rect 4786 14430 4820 14464
rect 4854 14430 4888 14464
rect 4922 14430 4956 14464
rect 4990 14430 5024 14464
rect 5058 14430 5092 14464
rect 5126 14430 5160 14464
rect 5194 14430 5228 14464
rect 5262 14430 5296 14464
rect 5330 14430 5364 14464
rect 5398 14430 5432 14464
rect 5466 14430 5500 14464
rect 5534 14430 5568 14464
rect 5602 14430 5636 14464
rect 5670 14430 5704 14464
rect 5738 14430 5772 14464
rect 5806 14430 5840 14464
rect 5874 14430 5908 14464
rect 5942 14430 5976 14464
rect 6010 14430 6044 14464
rect 6078 14430 6112 14464
rect 6146 14430 6180 14464
rect 6214 14430 6248 14464
rect 6282 14430 6316 14464
rect 6350 14430 6384 14464
rect 6418 14430 6452 14464
rect 6486 14430 6520 14464
rect 6554 14430 6588 14464
rect 6622 14430 6656 14464
rect 6690 14430 6724 14464
rect 6758 14430 6792 14464
rect 6826 14430 6860 14464
rect 6894 14430 6928 14464
rect 6962 14430 6996 14464
rect 7030 14430 7064 14464
rect 7098 14430 7132 14464
rect 7166 14430 7200 14464
rect 7234 14430 7268 14464
rect 7302 14430 7336 14464
rect 7370 14430 7404 14464
rect 7438 14430 7472 14464
rect 7506 14430 7540 14464
rect 7574 14430 7608 14464
rect 7642 14430 7676 14464
rect 7710 14430 7744 14464
rect 7778 14430 7812 14464
rect 7846 14430 7880 14464
rect 7914 14430 7948 14464
rect 7982 14430 8016 14464
rect 8050 14430 8084 14464
rect 8118 14430 8152 14464
rect 8186 14430 8220 14464
rect 8254 14430 8288 14464
rect 8322 14430 8356 14464
rect 8390 14430 8424 14464
rect 8458 14430 8492 14464
rect 8526 14430 8560 14464
rect 8594 14430 8628 14464
rect 8662 14430 8696 14464
rect 8730 14430 8764 14464
rect 8798 14430 8832 14464
rect 8866 14430 8900 14464
rect 8934 14430 8968 14464
rect 9002 14430 9036 14464
rect 9070 14430 9104 14464
rect 9138 14430 9172 14464
rect 9206 14430 9240 14464
rect 9274 14430 9308 14464
rect 9342 14430 9376 14464
rect 9410 14430 9444 14464
rect 9478 14430 9512 14464
rect 9546 14430 9580 14464
rect 9614 14430 9648 14464
rect 9682 14430 9716 14464
rect 9750 14430 9784 14464
rect 9818 14430 9852 14464
rect 9886 14430 9920 14464
rect 9954 14430 9988 14464
rect 10022 14430 10056 14464
rect 10090 14430 10124 14464
rect 10158 14430 10192 14464
rect 10226 14430 10260 14464
rect 10294 14430 10328 14464
rect 10362 14430 10396 14464
rect 10430 14430 10464 14464
rect 10498 14430 10532 14464
rect 10566 14430 10600 14464
rect 10634 14430 10668 14464
rect 10702 14430 10736 14464
rect 10770 14430 10804 14464
rect 10838 14430 10872 14464
rect 10906 14430 10940 14464
rect 10974 14430 11008 14464
rect 11042 14430 11076 14464
rect 11110 14430 11144 14464
rect 11178 14430 11212 14464
rect 11246 14430 11280 14464
rect 11314 14430 11348 14464
rect 11382 14430 11416 14464
rect 11450 14430 11484 14464
rect 11518 14430 11552 14464
rect 11586 14430 11620 14464
rect 11654 14430 11688 14464
rect 11722 14430 11756 14464
rect 11790 14430 11824 14464
rect 11858 14430 11892 14464
rect 11926 14430 11960 14464
rect 11994 14430 12028 14464
rect 12062 14430 12096 14464
rect 12130 14430 12164 14464
rect 12198 14430 12232 14464
rect 12266 14430 12300 14464
rect 12334 14430 12368 14464
rect 12402 14430 12436 14464
rect 12470 14430 12504 14464
rect 12538 14430 12572 14464
rect 12606 14430 12640 14464
rect 12674 14430 12708 14464
rect 12742 14430 12776 14464
rect 12810 14430 12844 14464
rect 12878 14430 12912 14464
rect 12946 14430 12980 14464
rect 13014 14430 13048 14464
rect 13082 14430 13116 14464
rect 13150 14430 13184 14464
rect 13218 14430 13252 14464
rect 13286 14430 13320 14464
rect 13354 14430 13388 14464
rect 13422 14430 13456 14464
rect 13490 14430 13524 14464
rect 13558 14430 13592 14464
rect 13626 14430 13660 14464
rect 13694 14430 13728 14464
rect 13762 14430 13796 14464
rect 13830 14430 13864 14464
rect 13898 14430 13932 14464
rect 13966 14430 14000 14464
rect 14034 14430 14068 14464
rect 14102 14430 14136 14464
rect 14170 14430 14204 14464
rect 14238 14430 14272 14464
rect 14306 14430 14340 14464
rect 14374 14430 14408 14464
rect 14442 14430 14476 14464
rect 14510 14430 14716 14464
rect 237 14356 14716 14430
<< mvnsubdiff >>
rect 575 36190 14373 36240
rect 575 36156 758 36190
rect 792 36156 826 36190
rect 860 36156 894 36190
rect 928 36156 962 36190
rect 996 36156 1030 36190
rect 1064 36156 1098 36190
rect 1132 36156 1166 36190
rect 1200 36156 1234 36190
rect 1268 36156 1302 36190
rect 1336 36156 1370 36190
rect 1404 36156 1438 36190
rect 1472 36156 1506 36190
rect 1540 36156 1574 36190
rect 1608 36156 1642 36190
rect 1676 36156 1710 36190
rect 1744 36156 1778 36190
rect 1812 36156 1846 36190
rect 1880 36156 1914 36190
rect 1948 36156 1982 36190
rect 2016 36156 2050 36190
rect 2084 36156 2118 36190
rect 2152 36156 2186 36190
rect 2220 36156 2254 36190
rect 2288 36156 2322 36190
rect 2356 36156 2390 36190
rect 2424 36156 2458 36190
rect 2492 36156 2526 36190
rect 2560 36156 2594 36190
rect 2628 36156 2662 36190
rect 2696 36156 2730 36190
rect 2764 36156 2798 36190
rect 2832 36156 2866 36190
rect 2900 36156 2934 36190
rect 2968 36156 3002 36190
rect 3036 36156 3070 36190
rect 3104 36156 3138 36190
rect 3172 36156 3206 36190
rect 3240 36156 3274 36190
rect 3308 36156 3342 36190
rect 3376 36156 3410 36190
rect 3444 36156 3478 36190
rect 3512 36156 3546 36190
rect 3580 36156 3614 36190
rect 3648 36156 3682 36190
rect 3716 36156 3750 36190
rect 3784 36156 3818 36190
rect 3852 36156 3886 36190
rect 3920 36156 3954 36190
rect 3988 36156 4022 36190
rect 4056 36156 4090 36190
rect 4124 36156 4158 36190
rect 4192 36156 4226 36190
rect 4260 36156 4294 36190
rect 4328 36156 4362 36190
rect 4396 36156 4430 36190
rect 4464 36156 4498 36190
rect 4532 36156 4566 36190
rect 4600 36156 4634 36190
rect 4668 36156 4702 36190
rect 4736 36156 4770 36190
rect 4804 36156 4838 36190
rect 4872 36156 4906 36190
rect 4940 36156 4974 36190
rect 5008 36156 5042 36190
rect 5076 36156 5110 36190
rect 5144 36156 5178 36190
rect 5212 36156 5246 36190
rect 5280 36156 5314 36190
rect 5348 36156 5382 36190
rect 5416 36156 5450 36190
rect 5484 36156 5518 36190
rect 5552 36156 5586 36190
rect 5620 36156 5654 36190
rect 5688 36156 5722 36190
rect 5756 36156 5790 36190
rect 5824 36156 5858 36190
rect 5892 36156 5926 36190
rect 5960 36156 5994 36190
rect 6028 36156 6062 36190
rect 6096 36156 6130 36190
rect 6164 36156 6198 36190
rect 6232 36156 6266 36190
rect 6300 36156 6334 36190
rect 6368 36156 6402 36190
rect 6436 36156 6470 36190
rect 6504 36156 6538 36190
rect 6572 36156 6606 36190
rect 6640 36156 6674 36190
rect 6708 36156 6742 36190
rect 6776 36156 6810 36190
rect 6844 36156 6878 36190
rect 6912 36156 6946 36190
rect 6980 36156 7014 36190
rect 7048 36156 7082 36190
rect 7116 36156 7150 36190
rect 7184 36156 7218 36190
rect 7252 36156 7286 36190
rect 7320 36156 7354 36190
rect 7388 36156 7422 36190
rect 7456 36156 7490 36190
rect 7524 36156 7558 36190
rect 7592 36156 7626 36190
rect 7660 36156 7694 36190
rect 7728 36156 7762 36190
rect 7796 36156 7830 36190
rect 7864 36156 7898 36190
rect 7932 36156 7966 36190
rect 8000 36156 8034 36190
rect 8068 36156 8102 36190
rect 8136 36156 8170 36190
rect 8204 36156 8238 36190
rect 8272 36156 8306 36190
rect 8340 36156 8374 36190
rect 8408 36156 8442 36190
rect 8476 36156 8510 36190
rect 8544 36156 8578 36190
rect 8612 36156 8646 36190
rect 8680 36156 8714 36190
rect 8748 36156 8782 36190
rect 8816 36156 8850 36190
rect 8884 36156 8918 36190
rect 8952 36156 8986 36190
rect 9020 36156 9054 36190
rect 9088 36156 9122 36190
rect 9156 36156 9190 36190
rect 9224 36156 9258 36190
rect 9292 36156 9326 36190
rect 9360 36156 9394 36190
rect 9428 36156 9462 36190
rect 9496 36156 9530 36190
rect 9564 36156 9598 36190
rect 9632 36156 9666 36190
rect 9700 36156 9734 36190
rect 9768 36156 9802 36190
rect 9836 36156 9870 36190
rect 9904 36156 9938 36190
rect 9972 36156 10006 36190
rect 10040 36156 10074 36190
rect 10108 36156 10142 36190
rect 10176 36156 10210 36190
rect 10244 36156 10278 36190
rect 10312 36156 10346 36190
rect 10380 36156 10414 36190
rect 10448 36156 10482 36190
rect 10516 36156 10550 36190
rect 10584 36156 10618 36190
rect 10652 36156 10686 36190
rect 10720 36156 10754 36190
rect 10788 36156 10822 36190
rect 10856 36156 10890 36190
rect 10924 36156 10958 36190
rect 10992 36156 11026 36190
rect 11060 36156 11094 36190
rect 11128 36156 11162 36190
rect 11196 36156 11230 36190
rect 11264 36156 11298 36190
rect 11332 36156 11366 36190
rect 11400 36156 11434 36190
rect 11468 36156 11502 36190
rect 11536 36156 11570 36190
rect 11604 36156 11638 36190
rect 11672 36156 11706 36190
rect 11740 36156 11774 36190
rect 11808 36156 11842 36190
rect 11876 36156 11910 36190
rect 11944 36156 11978 36190
rect 12012 36156 12046 36190
rect 12080 36156 12114 36190
rect 12148 36156 12182 36190
rect 12216 36156 12250 36190
rect 12284 36156 12318 36190
rect 12352 36156 12386 36190
rect 12420 36156 12454 36190
rect 12488 36156 12522 36190
rect 12556 36156 12590 36190
rect 12624 36156 12658 36190
rect 12692 36156 12726 36190
rect 12760 36156 12794 36190
rect 12828 36156 12862 36190
rect 12896 36156 12930 36190
rect 12964 36156 12998 36190
rect 13032 36156 13066 36190
rect 13100 36156 13134 36190
rect 13168 36156 13202 36190
rect 13236 36156 13270 36190
rect 13304 36156 13338 36190
rect 13372 36156 13406 36190
rect 13440 36156 13474 36190
rect 13508 36156 13542 36190
rect 13576 36156 13610 36190
rect 13644 36156 13678 36190
rect 13712 36156 13746 36190
rect 13780 36156 13814 36190
rect 13848 36156 13882 36190
rect 13916 36156 13950 36190
rect 13984 36156 14018 36190
rect 14052 36156 14086 36190
rect 14120 36156 14154 36190
rect 14188 36156 14373 36190
rect 575 36106 14373 36156
rect 575 36063 707 36106
rect 575 36029 624 36063
rect 658 36029 707 36063
rect 575 35995 707 36029
rect 575 35961 624 35995
rect 658 35961 707 35995
rect 575 35927 707 35961
rect 575 35893 624 35927
rect 658 35893 707 35927
rect 575 35859 707 35893
rect 575 35825 624 35859
rect 658 35825 707 35859
rect 575 35791 707 35825
rect 575 35757 624 35791
rect 658 35757 707 35791
rect 575 35723 707 35757
rect 575 35689 624 35723
rect 658 35689 707 35723
rect 575 35655 707 35689
rect 575 35621 624 35655
rect 658 35621 707 35655
rect 575 35587 707 35621
rect 575 35553 624 35587
rect 658 35553 707 35587
rect 575 35519 707 35553
rect 575 35485 624 35519
rect 658 35485 707 35519
rect 575 35451 707 35485
rect 575 35417 624 35451
rect 658 35417 707 35451
rect 575 35383 707 35417
rect 575 35349 624 35383
rect 658 35349 707 35383
rect 575 35315 707 35349
rect 575 35281 624 35315
rect 658 35281 707 35315
rect 575 35247 707 35281
rect 575 35213 624 35247
rect 658 35213 707 35247
rect 575 35179 707 35213
rect 575 35145 624 35179
rect 658 35145 707 35179
rect 575 35111 707 35145
rect 575 35077 624 35111
rect 658 35077 707 35111
rect 575 35043 707 35077
rect 575 35009 624 35043
rect 658 35009 707 35043
rect 575 34975 707 35009
rect 575 34941 624 34975
rect 658 34941 707 34975
rect 575 34907 707 34941
rect 575 34873 624 34907
rect 658 34873 707 34907
rect 575 34839 707 34873
rect 575 34805 624 34839
rect 658 34805 707 34839
rect 575 34771 707 34805
rect 575 34737 624 34771
rect 658 34737 707 34771
rect 575 34703 707 34737
rect 14239 36063 14373 36106
rect 14239 36029 14289 36063
rect 14323 36029 14373 36063
rect 14239 35995 14373 36029
rect 14239 35961 14289 35995
rect 14323 35961 14373 35995
rect 14239 35927 14373 35961
rect 14239 35893 14289 35927
rect 14323 35893 14373 35927
rect 14239 35859 14373 35893
rect 14239 35825 14289 35859
rect 14323 35825 14373 35859
rect 14239 35791 14373 35825
rect 14239 35757 14289 35791
rect 14323 35757 14373 35791
rect 14239 35723 14373 35757
rect 14239 35689 14289 35723
rect 14323 35689 14373 35723
rect 14239 35655 14373 35689
rect 14239 35621 14289 35655
rect 14323 35621 14373 35655
rect 14239 35587 14373 35621
rect 14239 35553 14289 35587
rect 14323 35553 14373 35587
rect 14239 35519 14373 35553
rect 14239 35485 14289 35519
rect 14323 35485 14373 35519
rect 14239 35451 14373 35485
rect 14239 35417 14289 35451
rect 14323 35417 14373 35451
rect 14239 35383 14373 35417
rect 14239 35349 14289 35383
rect 14323 35349 14373 35383
rect 14239 35315 14373 35349
rect 14239 35281 14289 35315
rect 14323 35281 14373 35315
rect 14239 35247 14373 35281
rect 14239 35213 14289 35247
rect 14323 35213 14373 35247
rect 14239 35179 14373 35213
rect 14239 35145 14289 35179
rect 14323 35145 14373 35179
rect 14239 35111 14373 35145
rect 14239 35077 14289 35111
rect 14323 35077 14373 35111
rect 14239 35043 14373 35077
rect 14239 35009 14289 35043
rect 14323 35009 14373 35043
rect 14239 34975 14373 35009
rect 14239 34941 14289 34975
rect 14323 34941 14373 34975
rect 14239 34907 14373 34941
rect 14239 34873 14289 34907
rect 14323 34873 14373 34907
rect 14239 34839 14373 34873
rect 14239 34805 14289 34839
rect 14323 34805 14373 34839
rect 14239 34771 14373 34805
rect 14239 34737 14289 34771
rect 14323 34737 14373 34771
rect 575 34669 624 34703
rect 658 34669 707 34703
rect 575 34635 707 34669
rect 575 34601 624 34635
rect 658 34601 707 34635
rect 575 34567 707 34601
rect 575 34533 624 34567
rect 658 34533 707 34567
rect 575 34499 707 34533
rect 575 34465 624 34499
rect 658 34465 707 34499
rect 575 34431 707 34465
rect 575 34397 624 34431
rect 658 34397 707 34431
rect 575 34363 707 34397
rect 575 34329 624 34363
rect 658 34329 707 34363
rect 575 34295 707 34329
rect 575 34261 624 34295
rect 658 34261 707 34295
rect 575 34227 707 34261
rect 575 34193 624 34227
rect 658 34193 707 34227
rect 575 34159 707 34193
rect 575 34125 624 34159
rect 658 34125 707 34159
rect 575 34091 707 34125
rect 575 34057 624 34091
rect 658 34057 707 34091
rect 575 34023 707 34057
rect 575 33989 624 34023
rect 658 33989 707 34023
rect 575 33955 707 33989
rect 575 33921 624 33955
rect 658 33921 707 33955
rect 575 33887 707 33921
rect 575 33853 624 33887
rect 658 33853 707 33887
rect 575 33819 707 33853
rect 575 33785 624 33819
rect 658 33785 707 33819
rect 575 33751 707 33785
rect 575 33717 624 33751
rect 658 33717 707 33751
rect 575 33683 707 33717
rect 575 33649 624 33683
rect 658 33649 707 33683
rect 575 33615 707 33649
rect 575 33581 624 33615
rect 658 33581 707 33615
rect 575 33547 707 33581
rect 575 33513 624 33547
rect 658 33513 707 33547
rect 575 33479 707 33513
rect 575 33445 624 33479
rect 658 33445 707 33479
rect 575 33411 707 33445
rect 575 33377 624 33411
rect 658 33377 707 33411
rect 575 33343 707 33377
rect 575 33309 624 33343
rect 658 33309 707 33343
rect 575 33275 707 33309
rect 575 33241 624 33275
rect 658 33241 707 33275
rect 575 33207 707 33241
rect 575 33173 624 33207
rect 658 33173 707 33207
rect 575 33139 707 33173
rect 575 33105 624 33139
rect 658 33105 707 33139
rect 575 33071 707 33105
rect 575 33037 624 33071
rect 658 33037 707 33071
rect 575 33003 707 33037
rect 575 32969 624 33003
rect 658 32969 707 33003
rect 575 32935 707 32969
rect 575 32901 624 32935
rect 658 32901 707 32935
rect 575 32867 707 32901
rect 575 32833 624 32867
rect 658 32833 707 32867
rect 575 32799 707 32833
rect 575 32765 624 32799
rect 658 32765 707 32799
rect 575 32731 707 32765
rect 575 32697 624 32731
rect 658 32697 707 32731
rect 575 32663 707 32697
rect 575 32629 624 32663
rect 658 32629 707 32663
rect 575 32595 707 32629
rect 575 32561 624 32595
rect 658 32561 707 32595
rect 575 32527 707 32561
rect 575 32493 624 32527
rect 658 32493 707 32527
rect 575 32459 707 32493
rect 575 32425 624 32459
rect 658 32425 707 32459
rect 575 32391 707 32425
rect 575 32357 624 32391
rect 658 32357 707 32391
rect 575 32323 707 32357
rect 575 32289 624 32323
rect 658 32289 707 32323
rect 575 32255 707 32289
rect 575 32221 624 32255
rect 658 32221 707 32255
rect 575 32187 707 32221
rect 575 32153 624 32187
rect 658 32153 707 32187
rect 575 32119 707 32153
rect 575 32085 624 32119
rect 658 32085 707 32119
rect 575 32051 707 32085
rect 575 32017 624 32051
rect 658 32017 707 32051
rect 575 31983 707 32017
rect 575 31949 624 31983
rect 658 31949 707 31983
rect 575 31915 707 31949
rect 575 31881 624 31915
rect 658 31881 707 31915
rect 575 31847 707 31881
rect 575 31813 624 31847
rect 658 31813 707 31847
rect 575 31779 707 31813
rect 575 31745 624 31779
rect 658 31745 707 31779
rect 575 31711 707 31745
rect 575 31677 624 31711
rect 658 31677 707 31711
rect 575 31643 707 31677
rect 575 31609 624 31643
rect 658 31609 707 31643
rect 575 31575 707 31609
rect 575 31541 624 31575
rect 658 31541 707 31575
rect 575 31507 707 31541
rect 575 31473 624 31507
rect 658 31473 707 31507
rect 575 31439 707 31473
rect 575 31405 624 31439
rect 658 31405 707 31439
rect 575 31371 707 31405
rect 575 31337 624 31371
rect 658 31337 707 31371
rect 575 31303 707 31337
rect 575 31269 624 31303
rect 658 31269 707 31303
rect 575 31235 707 31269
rect 575 31201 624 31235
rect 658 31201 707 31235
rect 575 31167 707 31201
rect 575 31133 624 31167
rect 658 31133 707 31167
rect 575 31099 707 31133
rect 575 31065 624 31099
rect 658 31065 707 31099
rect 575 31031 707 31065
rect 575 30997 624 31031
rect 658 30997 707 31031
rect 575 30963 707 30997
rect 575 30929 624 30963
rect 658 30929 707 30963
rect 575 30895 707 30929
rect 575 30861 624 30895
rect 658 30861 707 30895
rect 575 30827 707 30861
rect 575 30793 624 30827
rect 658 30793 707 30827
rect 575 30759 707 30793
rect 575 30725 624 30759
rect 658 30725 707 30759
rect 575 30691 707 30725
rect 575 30657 624 30691
rect 658 30657 707 30691
rect 575 30623 707 30657
rect 575 30589 624 30623
rect 658 30589 707 30623
rect 575 30555 707 30589
rect 575 30521 624 30555
rect 658 30521 707 30555
rect 575 30487 707 30521
rect 575 30453 624 30487
rect 658 30453 707 30487
rect 575 30419 707 30453
rect 575 30385 624 30419
rect 658 30385 707 30419
rect 575 30351 707 30385
rect 575 30317 624 30351
rect 658 30317 707 30351
rect 575 30283 707 30317
rect 575 30249 624 30283
rect 658 30249 707 30283
rect 575 30215 707 30249
rect 575 30181 624 30215
rect 658 30181 707 30215
rect 575 30147 707 30181
rect 575 30113 624 30147
rect 658 30113 707 30147
rect 575 30079 707 30113
rect 575 30045 624 30079
rect 658 30045 707 30079
rect 575 30011 707 30045
rect 575 29977 624 30011
rect 658 29977 707 30011
rect 575 29943 707 29977
rect 575 29909 624 29943
rect 658 29909 707 29943
rect 575 29875 707 29909
rect 575 29841 624 29875
rect 658 29841 707 29875
rect 575 29807 707 29841
rect 575 29773 624 29807
rect 658 29773 707 29807
rect 575 29739 707 29773
rect 575 29705 624 29739
rect 658 29705 707 29739
rect 575 29671 707 29705
rect 575 29637 624 29671
rect 658 29637 707 29671
rect 575 29603 707 29637
rect 575 29569 624 29603
rect 658 29569 707 29603
rect 575 29535 707 29569
rect 575 29501 624 29535
rect 658 29501 707 29535
rect 575 29467 707 29501
rect 575 29433 624 29467
rect 658 29433 707 29467
rect 575 29399 707 29433
rect 575 29365 624 29399
rect 658 29365 707 29399
rect 575 29331 707 29365
rect 575 29297 624 29331
rect 658 29297 707 29331
rect 575 29263 707 29297
rect 575 29229 624 29263
rect 658 29229 707 29263
rect 575 29195 707 29229
rect 575 29161 624 29195
rect 658 29161 707 29195
rect 575 29127 707 29161
rect 575 29093 624 29127
rect 658 29093 707 29127
rect 575 29059 707 29093
rect 575 29025 624 29059
rect 658 29025 707 29059
rect 575 28991 707 29025
rect 575 28957 624 28991
rect 658 28957 707 28991
rect 575 28923 707 28957
rect 575 28889 624 28923
rect 658 28889 707 28923
rect 575 28855 707 28889
rect 575 28821 624 28855
rect 658 28821 707 28855
rect 575 28787 707 28821
rect 575 28753 624 28787
rect 658 28753 707 28787
rect 575 28719 707 28753
rect 575 28685 624 28719
rect 658 28685 707 28719
rect 575 28651 707 28685
rect 575 28617 624 28651
rect 658 28617 707 28651
rect 575 28583 707 28617
rect 575 28549 624 28583
rect 658 28549 707 28583
rect 575 28515 707 28549
rect 575 28481 624 28515
rect 658 28481 707 28515
rect 575 28447 707 28481
rect 575 28413 624 28447
rect 658 28413 707 28447
rect 575 28379 707 28413
rect 575 28345 624 28379
rect 658 28345 707 28379
rect 575 28311 707 28345
rect 575 28277 624 28311
rect 658 28277 707 28311
rect 575 28243 707 28277
rect 575 28209 624 28243
rect 658 28209 707 28243
rect 575 28175 707 28209
rect 575 28141 624 28175
rect 658 28141 707 28175
rect 575 28107 707 28141
rect 575 28073 624 28107
rect 658 28073 707 28107
rect 575 28039 707 28073
rect 575 28005 624 28039
rect 658 28005 707 28039
rect 575 27971 707 28005
rect 575 27937 624 27971
rect 658 27937 707 27971
rect 575 27903 707 27937
rect 575 27869 624 27903
rect 658 27869 707 27903
rect 575 27835 707 27869
rect 575 27801 624 27835
rect 658 27801 707 27835
rect 575 27767 707 27801
rect 575 27733 624 27767
rect 658 27733 707 27767
rect 575 27699 707 27733
rect 575 27665 624 27699
rect 658 27665 707 27699
rect 575 27631 707 27665
rect 575 27597 624 27631
rect 658 27597 707 27631
rect 575 27563 707 27597
rect 575 27529 624 27563
rect 658 27529 707 27563
rect 575 27495 707 27529
rect 575 27461 624 27495
rect 658 27461 707 27495
rect 575 27427 707 27461
rect 575 27393 624 27427
rect 658 27393 707 27427
rect 575 27359 707 27393
rect 575 27325 624 27359
rect 658 27325 707 27359
rect 575 27291 707 27325
rect 575 27257 624 27291
rect 658 27257 707 27291
rect 575 27223 707 27257
rect 575 27189 624 27223
rect 658 27189 707 27223
rect 575 27155 707 27189
rect 575 27121 624 27155
rect 658 27121 707 27155
rect 575 27087 707 27121
rect 575 27053 624 27087
rect 658 27053 707 27087
rect 575 27019 707 27053
rect 575 26985 624 27019
rect 658 26985 707 27019
rect 575 26951 707 26985
rect 575 26917 624 26951
rect 658 26917 707 26951
rect 575 26883 707 26917
rect 575 26849 624 26883
rect 658 26849 707 26883
rect 575 26815 707 26849
rect 575 26781 624 26815
rect 658 26781 707 26815
rect 575 26747 707 26781
rect 575 26713 624 26747
rect 658 26713 707 26747
rect 575 26679 707 26713
rect 575 26645 624 26679
rect 658 26645 707 26679
rect 575 26611 707 26645
rect 575 26577 624 26611
rect 658 26577 707 26611
rect 575 26543 707 26577
rect 575 26509 624 26543
rect 658 26509 707 26543
rect 575 26475 707 26509
rect 575 26441 624 26475
rect 658 26441 707 26475
rect 575 26407 707 26441
rect 575 26373 624 26407
rect 658 26373 707 26407
rect 575 26339 707 26373
rect 575 26305 624 26339
rect 658 26305 707 26339
rect 575 26271 707 26305
rect 575 26237 624 26271
rect 658 26237 707 26271
rect 575 26203 707 26237
rect 575 26169 624 26203
rect 658 26169 707 26203
rect 575 26135 707 26169
rect 575 26101 624 26135
rect 658 26101 707 26135
rect 575 26067 707 26101
rect 575 26033 624 26067
rect 658 26033 707 26067
rect 575 25999 707 26033
rect 575 25965 624 25999
rect 658 25965 707 25999
rect 575 25931 707 25965
rect 575 25897 624 25931
rect 658 25897 707 25931
rect 575 25863 707 25897
rect 575 25829 624 25863
rect 658 25829 707 25863
rect 575 25795 707 25829
rect 575 25761 624 25795
rect 658 25761 707 25795
rect 575 25727 707 25761
rect 575 25693 624 25727
rect 658 25693 707 25727
rect 575 25659 707 25693
rect 575 25625 624 25659
rect 658 25625 707 25659
rect 575 25591 707 25625
rect 575 25557 624 25591
rect 658 25557 707 25591
rect 575 25523 707 25557
rect 575 25489 624 25523
rect 658 25489 707 25523
rect 575 25455 707 25489
rect 575 25421 624 25455
rect 658 25421 707 25455
rect 575 25387 707 25421
rect 575 25353 624 25387
rect 658 25353 707 25387
rect 575 25319 707 25353
rect 575 25285 624 25319
rect 658 25285 707 25319
rect 575 25251 707 25285
rect 575 25217 624 25251
rect 658 25217 707 25251
rect 575 25183 707 25217
rect 575 25149 624 25183
rect 658 25149 707 25183
rect 575 25115 707 25149
rect 575 25081 624 25115
rect 658 25081 707 25115
rect 575 25047 707 25081
rect 575 25013 624 25047
rect 658 25013 707 25047
rect 575 24979 707 25013
rect 575 24945 624 24979
rect 658 24945 707 24979
rect 575 24911 707 24945
rect 575 24877 624 24911
rect 658 24877 707 24911
rect 575 24843 707 24877
rect 575 24809 624 24843
rect 658 24809 707 24843
rect 575 24775 707 24809
rect 575 24741 624 24775
rect 658 24741 707 24775
rect 575 24707 707 24741
rect 575 24673 624 24707
rect 658 24673 707 24707
rect 575 24639 707 24673
rect 575 24605 624 24639
rect 658 24605 707 24639
rect 575 24571 707 24605
rect 575 24537 624 24571
rect 658 24537 707 24571
rect 575 24503 707 24537
rect 575 24469 624 24503
rect 658 24469 707 24503
rect 575 24435 707 24469
rect 575 24401 624 24435
rect 658 24401 707 24435
rect 575 24367 707 24401
rect 575 24333 624 24367
rect 658 24333 707 24367
rect 575 24299 707 24333
rect 575 24265 624 24299
rect 658 24265 707 24299
rect 575 24231 707 24265
rect 575 24197 624 24231
rect 658 24197 707 24231
rect 575 24163 707 24197
rect 575 24129 624 24163
rect 658 24129 707 24163
rect 575 24095 707 24129
rect 575 24061 624 24095
rect 658 24061 707 24095
rect 575 24027 707 24061
rect 575 23993 624 24027
rect 658 23993 707 24027
rect 575 23959 707 23993
rect 575 23925 624 23959
rect 658 23925 707 23959
rect 575 23891 707 23925
rect 575 23857 624 23891
rect 658 23857 707 23891
rect 575 23823 707 23857
rect 575 23789 624 23823
rect 658 23789 707 23823
rect 575 23755 707 23789
rect 575 23721 624 23755
rect 658 23721 707 23755
rect 575 23687 707 23721
rect 575 23653 624 23687
rect 658 23653 707 23687
rect 575 23619 707 23653
rect 575 23585 624 23619
rect 658 23585 707 23619
rect 575 23551 707 23585
rect 575 23517 624 23551
rect 658 23517 707 23551
rect 575 23483 707 23517
rect 575 23449 624 23483
rect 658 23449 707 23483
rect 575 23415 707 23449
rect 575 23381 624 23415
rect 658 23381 707 23415
rect 575 23347 707 23381
rect 575 23313 624 23347
rect 658 23313 707 23347
rect 575 23279 707 23313
rect 575 23245 624 23279
rect 658 23245 707 23279
rect 575 23211 707 23245
rect 575 23177 624 23211
rect 658 23177 707 23211
rect 575 23143 707 23177
rect 575 23109 624 23143
rect 658 23109 707 23143
rect 575 23075 707 23109
rect 575 23041 624 23075
rect 658 23041 707 23075
rect 575 23007 707 23041
rect 575 22973 624 23007
rect 658 22973 707 23007
rect 575 22939 707 22973
rect 575 22905 624 22939
rect 658 22905 707 22939
rect 575 22871 707 22905
rect 575 22837 624 22871
rect 658 22837 707 22871
rect 575 22803 707 22837
rect 575 22769 624 22803
rect 658 22769 707 22803
rect 575 22735 707 22769
rect 575 22701 624 22735
rect 658 22701 707 22735
rect 575 22667 707 22701
rect 575 22633 624 22667
rect 658 22633 707 22667
rect 575 22599 707 22633
rect 575 22565 624 22599
rect 658 22565 707 22599
rect 575 22531 707 22565
rect 575 22497 624 22531
rect 658 22497 707 22531
rect 575 22463 707 22497
rect 575 22429 624 22463
rect 658 22429 707 22463
rect 575 22395 707 22429
rect 575 22361 624 22395
rect 658 22361 707 22395
rect 575 22327 707 22361
rect 575 22293 624 22327
rect 658 22293 707 22327
rect 575 22259 707 22293
rect 575 22225 624 22259
rect 658 22225 707 22259
rect 575 22191 707 22225
rect 575 22157 624 22191
rect 658 22157 707 22191
rect 575 22123 707 22157
rect 575 22089 624 22123
rect 658 22089 707 22123
rect 575 22055 707 22089
rect 575 22021 624 22055
rect 658 22021 707 22055
rect 575 21987 707 22021
rect 575 21953 624 21987
rect 658 21953 707 21987
rect 575 21919 707 21953
rect 575 21885 624 21919
rect 658 21885 707 21919
rect 575 21851 707 21885
rect 575 21817 624 21851
rect 658 21817 707 21851
rect 575 21783 707 21817
rect 575 21749 624 21783
rect 658 21749 707 21783
rect 575 21715 707 21749
rect 575 21681 624 21715
rect 658 21681 707 21715
rect 575 21647 707 21681
rect 575 21613 624 21647
rect 658 21613 707 21647
rect 575 21579 707 21613
rect 575 21545 624 21579
rect 658 21545 707 21579
rect 575 21511 707 21545
rect 575 21477 624 21511
rect 658 21477 707 21511
rect 575 21443 707 21477
rect 575 21409 624 21443
rect 658 21409 707 21443
rect 575 21375 707 21409
rect 575 21341 624 21375
rect 658 21341 707 21375
rect 575 21307 707 21341
rect 575 21273 624 21307
rect 658 21273 707 21307
rect 575 21239 707 21273
rect 575 21205 624 21239
rect 658 21205 707 21239
rect 575 21171 707 21205
rect 575 21137 624 21171
rect 658 21137 707 21171
rect 575 21103 707 21137
rect 575 21069 624 21103
rect 658 21069 707 21103
rect 575 21035 707 21069
rect 575 21001 624 21035
rect 658 21001 707 21035
rect 575 20967 707 21001
rect 575 20933 624 20967
rect 658 20933 707 20967
rect 575 20899 707 20933
rect 575 20865 624 20899
rect 658 20865 707 20899
rect 575 20831 707 20865
rect 575 20797 624 20831
rect 658 20797 707 20831
rect 575 20763 707 20797
rect 575 20729 624 20763
rect 658 20729 707 20763
rect 575 20695 707 20729
rect 575 20661 624 20695
rect 658 20661 707 20695
rect 575 20627 707 20661
rect 575 20593 624 20627
rect 658 20593 707 20627
rect 575 20559 707 20593
rect 575 20525 624 20559
rect 658 20525 707 20559
rect 575 20491 707 20525
rect 575 20457 624 20491
rect 658 20457 707 20491
rect 575 20423 707 20457
rect 575 20389 624 20423
rect 658 20389 707 20423
rect 575 20355 707 20389
rect 575 20321 624 20355
rect 658 20321 707 20355
rect 575 20287 707 20321
rect 575 20253 624 20287
rect 658 20253 707 20287
rect 575 20219 707 20253
rect 575 20185 624 20219
rect 658 20185 707 20219
rect 575 20151 707 20185
rect 575 20117 624 20151
rect 658 20117 707 20151
rect 575 20083 707 20117
rect 575 20049 624 20083
rect 658 20049 707 20083
rect 575 20015 707 20049
rect 575 19981 624 20015
rect 658 19981 707 20015
rect 575 19947 707 19981
rect 575 19913 624 19947
rect 658 19913 707 19947
rect 575 19879 707 19913
rect 575 19845 624 19879
rect 658 19845 707 19879
rect 575 19811 707 19845
rect 575 19777 624 19811
rect 658 19777 707 19811
rect 575 19743 707 19777
rect 575 19709 624 19743
rect 658 19709 707 19743
rect 575 19675 707 19709
rect 575 19641 624 19675
rect 658 19641 707 19675
rect 575 19607 707 19641
rect 575 19573 624 19607
rect 658 19573 707 19607
rect 575 19539 707 19573
rect 575 19505 624 19539
rect 658 19505 707 19539
rect 575 19471 707 19505
rect 575 19437 624 19471
rect 658 19437 707 19471
rect 575 19403 707 19437
rect 575 19369 624 19403
rect 658 19369 707 19403
rect 575 19335 707 19369
rect 575 19301 624 19335
rect 658 19301 707 19335
rect 575 19267 707 19301
rect 575 19233 624 19267
rect 658 19233 707 19267
rect 575 19199 707 19233
rect 575 19165 624 19199
rect 658 19165 707 19199
rect 575 19131 707 19165
rect 575 19097 624 19131
rect 658 19097 707 19131
rect 575 19063 707 19097
rect 575 19029 624 19063
rect 658 19029 707 19063
rect 575 18995 707 19029
rect 575 18961 624 18995
rect 658 18961 707 18995
rect 575 18927 707 18961
rect 575 18893 624 18927
rect 658 18893 707 18927
rect 575 18859 707 18893
rect 575 18825 624 18859
rect 658 18825 707 18859
rect 575 18791 707 18825
rect 575 18757 624 18791
rect 658 18757 707 18791
rect 575 18723 707 18757
rect 575 18689 624 18723
rect 658 18689 707 18723
rect 575 18655 707 18689
rect 575 18621 624 18655
rect 658 18621 707 18655
rect 575 18587 707 18621
rect 575 18553 624 18587
rect 658 18553 707 18587
rect 575 18519 707 18553
rect 575 18485 624 18519
rect 658 18485 707 18519
rect 575 18451 707 18485
rect 575 18417 624 18451
rect 658 18417 707 18451
rect 575 18383 707 18417
rect 575 18349 624 18383
rect 658 18349 707 18383
rect 575 18315 707 18349
rect 575 18281 624 18315
rect 658 18281 707 18315
rect 575 18247 707 18281
rect 575 18213 624 18247
rect 658 18213 707 18247
rect 575 18179 707 18213
rect 575 18145 624 18179
rect 658 18145 707 18179
rect 575 18111 707 18145
rect 575 18077 624 18111
rect 658 18077 707 18111
rect 575 18043 707 18077
rect 575 18009 624 18043
rect 658 18009 707 18043
rect 575 17975 707 18009
rect 575 17941 624 17975
rect 658 17941 707 17975
rect 575 17907 707 17941
rect 575 17873 624 17907
rect 658 17873 707 17907
rect 575 17839 707 17873
rect 575 17805 624 17839
rect 658 17805 707 17839
rect 575 17771 707 17805
rect 575 17737 624 17771
rect 658 17737 707 17771
rect 575 17703 707 17737
rect 575 17669 624 17703
rect 658 17669 707 17703
rect 575 17635 707 17669
rect 575 17601 624 17635
rect 658 17601 707 17635
rect 575 17567 707 17601
rect 575 17533 624 17567
rect 658 17533 707 17567
rect 575 17499 707 17533
rect 575 17465 624 17499
rect 658 17465 707 17499
rect 575 17431 707 17465
rect 575 17397 624 17431
rect 658 17397 707 17431
rect 575 17363 707 17397
rect 575 17329 624 17363
rect 658 17329 707 17363
rect 575 17295 707 17329
rect 575 17261 624 17295
rect 658 17261 707 17295
rect 575 17227 707 17261
rect 575 17193 624 17227
rect 658 17193 707 17227
rect 575 17159 707 17193
rect 575 17125 624 17159
rect 658 17125 707 17159
rect 575 17091 707 17125
rect 575 17057 624 17091
rect 658 17057 707 17091
rect 575 17023 707 17057
rect 575 16989 624 17023
rect 658 16989 707 17023
rect 575 16955 707 16989
rect 575 16921 624 16955
rect 658 16921 707 16955
rect 575 16887 707 16921
rect 575 16853 624 16887
rect 658 16853 707 16887
rect 575 16819 707 16853
rect 575 16785 624 16819
rect 658 16785 707 16819
rect 575 16751 707 16785
rect 575 16717 624 16751
rect 658 16717 707 16751
rect 575 16683 707 16717
rect 575 16649 624 16683
rect 658 16649 707 16683
rect 575 16615 707 16649
rect 575 16581 624 16615
rect 658 16581 707 16615
rect 575 16547 707 16581
rect 575 16513 624 16547
rect 658 16513 707 16547
rect 575 16479 707 16513
rect 575 16445 624 16479
rect 658 16445 707 16479
rect 575 16411 707 16445
rect 575 16377 624 16411
rect 658 16377 707 16411
rect 575 16343 707 16377
rect 575 16309 624 16343
rect 658 16309 707 16343
rect 575 16275 707 16309
rect 575 16241 624 16275
rect 658 16241 707 16275
rect 575 16207 707 16241
rect 575 16173 624 16207
rect 658 16173 707 16207
rect 575 16139 707 16173
rect 575 16105 624 16139
rect 658 16105 707 16139
rect 575 16071 707 16105
rect 575 16037 624 16071
rect 658 16037 707 16071
rect 575 16003 707 16037
rect 575 15969 624 16003
rect 658 15969 707 16003
rect 575 15935 707 15969
rect 575 15901 624 15935
rect 658 15901 707 15935
rect 575 15867 707 15901
rect 575 15833 624 15867
rect 658 15833 707 15867
rect 575 15799 707 15833
rect 575 15765 624 15799
rect 658 15765 707 15799
rect 575 15731 707 15765
rect 575 15697 624 15731
rect 658 15697 707 15731
rect 575 15663 707 15697
rect 575 15629 624 15663
rect 658 15629 707 15663
rect 575 15595 707 15629
rect 575 15561 624 15595
rect 658 15561 707 15595
rect 575 15527 707 15561
rect 575 15493 624 15527
rect 658 15493 707 15527
rect 575 15459 707 15493
rect 575 15425 624 15459
rect 658 15425 707 15459
rect 575 15391 707 15425
rect 575 15357 624 15391
rect 658 15357 707 15391
rect 575 15323 707 15357
rect 575 15289 624 15323
rect 658 15289 707 15323
rect 575 15255 707 15289
rect 575 15221 624 15255
rect 658 15221 707 15255
rect 575 15187 707 15221
rect 1651 28892 13349 28922
rect 1651 28518 2111 28892
rect 12889 28518 13349 28892
rect 1651 28488 13349 28518
rect 1651 28435 2085 28488
rect 1651 27517 1681 28435
rect 2055 27517 2085 28435
rect 12915 28435 13349 28488
rect 1651 27464 2085 27517
rect 12915 27517 12945 28435
rect 13319 27517 13349 28435
rect 12915 27464 13349 27517
rect 1651 27434 13349 27464
rect 1651 27060 2111 27434
rect 12889 27060 13349 27434
rect 1651 27030 13349 27060
rect 2386 25909 12590 25979
rect 2386 25875 2473 25909
rect 2507 25875 2541 25909
rect 2575 25875 2609 25909
rect 2643 25875 2677 25909
rect 2711 25875 2745 25909
rect 2779 25875 2813 25909
rect 2847 25875 2881 25909
rect 2915 25875 2949 25909
rect 2983 25875 3017 25909
rect 3051 25875 3085 25909
rect 3119 25875 3153 25909
rect 3187 25875 3221 25909
rect 3255 25875 3289 25909
rect 3323 25875 3357 25909
rect 3391 25875 3425 25909
rect 3459 25875 3493 25909
rect 3527 25875 3561 25909
rect 3595 25875 3629 25909
rect 3663 25875 3697 25909
rect 3731 25875 3765 25909
rect 3799 25875 3833 25909
rect 3867 25875 3901 25909
rect 3935 25875 3969 25909
rect 4003 25875 4037 25909
rect 4071 25875 4105 25909
rect 4139 25875 4173 25909
rect 4207 25875 4241 25909
rect 4275 25875 4309 25909
rect 4343 25875 4377 25909
rect 4411 25875 4445 25909
rect 4479 25875 4513 25909
rect 4547 25875 4581 25909
rect 4615 25875 4649 25909
rect 4683 25875 4717 25909
rect 4751 25875 4785 25909
rect 4819 25875 4853 25909
rect 4887 25875 4921 25909
rect 4955 25875 4989 25909
rect 5023 25875 5057 25909
rect 5091 25875 5125 25909
rect 5159 25875 5193 25909
rect 5227 25875 5261 25909
rect 5295 25875 5329 25909
rect 5363 25875 5397 25909
rect 5431 25875 5465 25909
rect 5499 25875 5533 25909
rect 5567 25875 5601 25909
rect 5635 25875 5669 25909
rect 5703 25875 5737 25909
rect 5771 25875 5805 25909
rect 5839 25875 5873 25909
rect 5907 25875 5941 25909
rect 5975 25875 6009 25909
rect 6043 25875 6077 25909
rect 6111 25875 6145 25909
rect 6179 25875 6213 25909
rect 6247 25875 6281 25909
rect 6315 25875 6349 25909
rect 6383 25875 6417 25909
rect 6451 25875 6485 25909
rect 6519 25875 6553 25909
rect 6587 25875 6621 25909
rect 6655 25875 6689 25909
rect 6723 25875 6757 25909
rect 6791 25875 6825 25909
rect 6859 25875 6893 25909
rect 6927 25875 6961 25909
rect 6995 25875 7029 25909
rect 7063 25875 7097 25909
rect 7131 25875 7165 25909
rect 7199 25875 7233 25909
rect 7267 25875 7301 25909
rect 7335 25875 7369 25909
rect 7403 25875 7437 25909
rect 7471 25875 7505 25909
rect 7539 25875 7573 25909
rect 7607 25875 7641 25909
rect 7675 25875 7709 25909
rect 7743 25875 7777 25909
rect 7811 25875 7845 25909
rect 7879 25875 7913 25909
rect 7947 25875 7981 25909
rect 8015 25875 8049 25909
rect 8083 25875 8117 25909
rect 8151 25875 8185 25909
rect 8219 25875 8253 25909
rect 8287 25875 8321 25909
rect 8355 25875 8389 25909
rect 8423 25875 8457 25909
rect 8491 25875 8525 25909
rect 8559 25875 8593 25909
rect 8627 25875 8661 25909
rect 8695 25875 8729 25909
rect 8763 25875 8797 25909
rect 8831 25875 8865 25909
rect 8899 25875 8933 25909
rect 8967 25875 9001 25909
rect 9035 25875 9069 25909
rect 9103 25875 9137 25909
rect 9171 25875 9205 25909
rect 9239 25875 9273 25909
rect 9307 25875 9341 25909
rect 9375 25875 9409 25909
rect 9443 25875 9477 25909
rect 9511 25875 9545 25909
rect 9579 25875 9613 25909
rect 9647 25875 9681 25909
rect 9715 25875 9749 25909
rect 9783 25875 9817 25909
rect 9851 25875 9885 25909
rect 9919 25875 9953 25909
rect 9987 25875 10021 25909
rect 10055 25875 10089 25909
rect 10123 25875 10157 25909
rect 10191 25875 10225 25909
rect 10259 25875 10293 25909
rect 10327 25875 10361 25909
rect 10395 25875 10429 25909
rect 10463 25875 10497 25909
rect 10531 25875 10565 25909
rect 10599 25875 10633 25909
rect 10667 25875 10701 25909
rect 10735 25875 10769 25909
rect 10803 25875 10837 25909
rect 10871 25875 10905 25909
rect 10939 25875 10973 25909
rect 11007 25875 11041 25909
rect 11075 25875 11109 25909
rect 11143 25875 11177 25909
rect 11211 25875 11245 25909
rect 11279 25875 11313 25909
rect 11347 25875 11381 25909
rect 11415 25875 11449 25909
rect 11483 25875 11517 25909
rect 11551 25875 11585 25909
rect 11619 25875 11653 25909
rect 11687 25875 11721 25909
rect 11755 25875 11789 25909
rect 11823 25875 11857 25909
rect 11891 25875 11925 25909
rect 11959 25875 11993 25909
rect 12027 25875 12061 25909
rect 12095 25875 12129 25909
rect 12163 25875 12197 25909
rect 12231 25875 12265 25909
rect 12299 25875 12333 25909
rect 12367 25875 12401 25909
rect 12435 25875 12469 25909
rect 12503 25875 12590 25909
rect 2386 25826 2420 25875
rect 12556 25826 12590 25875
rect 2386 25758 2420 25792
rect 2386 25690 2420 25724
rect 2386 25622 2420 25656
rect 12556 25758 12590 25792
rect 12556 25690 12590 25724
rect 12556 25622 12590 25656
rect 2386 25539 2420 25588
rect 12556 25539 12590 25588
rect 2386 25505 2473 25539
rect 2507 25505 2541 25539
rect 2575 25505 2609 25539
rect 2643 25505 2677 25539
rect 2711 25505 2745 25539
rect 2779 25505 2813 25539
rect 2847 25505 2881 25539
rect 2915 25505 2949 25539
rect 2983 25505 3017 25539
rect 3051 25505 3085 25539
rect 3119 25505 3153 25539
rect 3187 25505 3221 25539
rect 3255 25505 3289 25539
rect 3323 25505 3357 25539
rect 3391 25505 3425 25539
rect 3459 25505 3493 25539
rect 3527 25505 3561 25539
rect 3595 25505 3629 25539
rect 3663 25505 3697 25539
rect 3731 25505 3765 25539
rect 3799 25505 3833 25539
rect 3867 25505 3901 25539
rect 3935 25505 3969 25539
rect 4003 25505 4037 25539
rect 4071 25505 4105 25539
rect 4139 25505 4173 25539
rect 4207 25505 4241 25539
rect 4275 25505 4309 25539
rect 4343 25505 4377 25539
rect 4411 25505 4445 25539
rect 4479 25505 4513 25539
rect 4547 25505 4581 25539
rect 4615 25505 4649 25539
rect 4683 25505 4717 25539
rect 4751 25505 4785 25539
rect 4819 25505 4853 25539
rect 4887 25505 4921 25539
rect 4955 25505 4989 25539
rect 5023 25505 5057 25539
rect 5091 25505 5125 25539
rect 5159 25505 5193 25539
rect 5227 25505 5261 25539
rect 5295 25505 5329 25539
rect 5363 25505 5397 25539
rect 5431 25505 5465 25539
rect 5499 25505 5533 25539
rect 5567 25505 5601 25539
rect 5635 25505 5669 25539
rect 5703 25505 5737 25539
rect 5771 25505 5805 25539
rect 5839 25505 5873 25539
rect 5907 25505 5941 25539
rect 5975 25505 6009 25539
rect 6043 25505 6077 25539
rect 6111 25505 6145 25539
rect 6179 25505 6213 25539
rect 6247 25505 6281 25539
rect 6315 25505 6349 25539
rect 6383 25505 6417 25539
rect 6451 25505 6485 25539
rect 6519 25505 6553 25539
rect 6587 25505 6621 25539
rect 6655 25505 6689 25539
rect 6723 25505 6757 25539
rect 6791 25505 6825 25539
rect 6859 25505 6893 25539
rect 6927 25505 6961 25539
rect 6995 25505 7029 25539
rect 7063 25505 7097 25539
rect 7131 25505 7165 25539
rect 7199 25505 7233 25539
rect 7267 25505 7301 25539
rect 7335 25505 7369 25539
rect 7403 25505 7437 25539
rect 7471 25505 7505 25539
rect 7539 25505 7573 25539
rect 7607 25505 7641 25539
rect 7675 25505 7709 25539
rect 7743 25505 7777 25539
rect 7811 25505 7845 25539
rect 7879 25505 7913 25539
rect 7947 25505 7981 25539
rect 8015 25505 8049 25539
rect 8083 25505 8117 25539
rect 8151 25505 8185 25539
rect 8219 25505 8253 25539
rect 8287 25505 8321 25539
rect 8355 25505 8389 25539
rect 8423 25505 8457 25539
rect 8491 25505 8525 25539
rect 8559 25505 8593 25539
rect 8627 25505 8661 25539
rect 8695 25505 8729 25539
rect 8763 25505 8797 25539
rect 8831 25505 8865 25539
rect 8899 25505 8933 25539
rect 8967 25505 9001 25539
rect 9035 25505 9069 25539
rect 9103 25505 9137 25539
rect 9171 25505 9205 25539
rect 9239 25505 9273 25539
rect 9307 25505 9341 25539
rect 9375 25505 9409 25539
rect 9443 25505 9477 25539
rect 9511 25505 9545 25539
rect 9579 25505 9613 25539
rect 9647 25505 9681 25539
rect 9715 25505 9749 25539
rect 9783 25505 9817 25539
rect 9851 25505 9885 25539
rect 9919 25505 9953 25539
rect 9987 25505 10021 25539
rect 10055 25505 10089 25539
rect 10123 25505 10157 25539
rect 10191 25505 10225 25539
rect 10259 25505 10293 25539
rect 10327 25505 10361 25539
rect 10395 25505 10429 25539
rect 10463 25505 10497 25539
rect 10531 25505 10565 25539
rect 10599 25505 10633 25539
rect 10667 25505 10701 25539
rect 10735 25505 10769 25539
rect 10803 25505 10837 25539
rect 10871 25505 10905 25539
rect 10939 25505 10973 25539
rect 11007 25505 11041 25539
rect 11075 25505 11109 25539
rect 11143 25505 11177 25539
rect 11211 25505 11245 25539
rect 11279 25505 11313 25539
rect 11347 25505 11381 25539
rect 11415 25505 11449 25539
rect 11483 25505 11517 25539
rect 11551 25505 11585 25539
rect 11619 25505 11653 25539
rect 11687 25505 11721 25539
rect 11755 25505 11789 25539
rect 11823 25505 11857 25539
rect 11891 25505 11925 25539
rect 11959 25505 11993 25539
rect 12027 25505 12061 25539
rect 12095 25505 12129 25539
rect 12163 25505 12197 25539
rect 12231 25505 12265 25539
rect 12299 25505 12333 25539
rect 12367 25505 12401 25539
rect 12435 25505 12469 25539
rect 12503 25505 12590 25539
rect 2386 25441 12590 25505
rect 14239 34703 14373 34737
rect 14239 34669 14289 34703
rect 14323 34669 14373 34703
rect 14239 34635 14373 34669
rect 14239 34601 14289 34635
rect 14323 34601 14373 34635
rect 14239 34567 14373 34601
rect 14239 34533 14289 34567
rect 14323 34533 14373 34567
rect 14239 34499 14373 34533
rect 14239 34465 14289 34499
rect 14323 34465 14373 34499
rect 14239 34431 14373 34465
rect 14239 34397 14289 34431
rect 14323 34397 14373 34431
rect 14239 34363 14373 34397
rect 14239 34329 14289 34363
rect 14323 34329 14373 34363
rect 14239 34295 14373 34329
rect 14239 34261 14289 34295
rect 14323 34261 14373 34295
rect 14239 34227 14373 34261
rect 14239 34193 14289 34227
rect 14323 34193 14373 34227
rect 14239 34159 14373 34193
rect 14239 34125 14289 34159
rect 14323 34125 14373 34159
rect 14239 34091 14373 34125
rect 14239 34057 14289 34091
rect 14323 34057 14373 34091
rect 14239 34023 14373 34057
rect 14239 33989 14289 34023
rect 14323 33989 14373 34023
rect 14239 33955 14373 33989
rect 14239 33921 14289 33955
rect 14323 33921 14373 33955
rect 14239 33887 14373 33921
rect 14239 33853 14289 33887
rect 14323 33853 14373 33887
rect 14239 33819 14373 33853
rect 14239 33785 14289 33819
rect 14323 33785 14373 33819
rect 14239 33751 14373 33785
rect 14239 33717 14289 33751
rect 14323 33717 14373 33751
rect 14239 33683 14373 33717
rect 14239 33649 14289 33683
rect 14323 33649 14373 33683
rect 14239 33615 14373 33649
rect 14239 33581 14289 33615
rect 14323 33581 14373 33615
rect 14239 33547 14373 33581
rect 14239 33513 14289 33547
rect 14323 33513 14373 33547
rect 14239 33479 14373 33513
rect 14239 33445 14289 33479
rect 14323 33445 14373 33479
rect 14239 33411 14373 33445
rect 14239 33377 14289 33411
rect 14323 33377 14373 33411
rect 14239 33343 14373 33377
rect 14239 33309 14289 33343
rect 14323 33309 14373 33343
rect 14239 33275 14373 33309
rect 14239 33241 14289 33275
rect 14323 33241 14373 33275
rect 14239 33207 14373 33241
rect 14239 33173 14289 33207
rect 14323 33173 14373 33207
rect 14239 33139 14373 33173
rect 14239 33105 14289 33139
rect 14323 33105 14373 33139
rect 14239 33071 14373 33105
rect 14239 33037 14289 33071
rect 14323 33037 14373 33071
rect 14239 33003 14373 33037
rect 14239 32969 14289 33003
rect 14323 32969 14373 33003
rect 14239 32935 14373 32969
rect 14239 32901 14289 32935
rect 14323 32901 14373 32935
rect 14239 32867 14373 32901
rect 14239 32833 14289 32867
rect 14323 32833 14373 32867
rect 14239 32799 14373 32833
rect 14239 32765 14289 32799
rect 14323 32765 14373 32799
rect 14239 32731 14373 32765
rect 14239 32697 14289 32731
rect 14323 32697 14373 32731
rect 14239 32663 14373 32697
rect 14239 32629 14289 32663
rect 14323 32629 14373 32663
rect 14239 32595 14373 32629
rect 14239 32561 14289 32595
rect 14323 32561 14373 32595
rect 14239 32527 14373 32561
rect 14239 32493 14289 32527
rect 14323 32493 14373 32527
rect 14239 32459 14373 32493
rect 14239 32425 14289 32459
rect 14323 32425 14373 32459
rect 14239 32391 14373 32425
rect 14239 32357 14289 32391
rect 14323 32357 14373 32391
rect 14239 32323 14373 32357
rect 14239 32289 14289 32323
rect 14323 32289 14373 32323
rect 14239 32255 14373 32289
rect 14239 32221 14289 32255
rect 14323 32221 14373 32255
rect 14239 32187 14373 32221
rect 14239 32153 14289 32187
rect 14323 32153 14373 32187
rect 14239 32119 14373 32153
rect 14239 32085 14289 32119
rect 14323 32085 14373 32119
rect 14239 32051 14373 32085
rect 14239 32017 14289 32051
rect 14323 32017 14373 32051
rect 14239 31983 14373 32017
rect 14239 31949 14289 31983
rect 14323 31949 14373 31983
rect 14239 31915 14373 31949
rect 14239 31881 14289 31915
rect 14323 31881 14373 31915
rect 14239 31847 14373 31881
rect 14239 31813 14289 31847
rect 14323 31813 14373 31847
rect 14239 31779 14373 31813
rect 14239 31745 14289 31779
rect 14323 31745 14373 31779
rect 14239 31711 14373 31745
rect 14239 31677 14289 31711
rect 14323 31677 14373 31711
rect 14239 31643 14373 31677
rect 14239 31609 14289 31643
rect 14323 31609 14373 31643
rect 14239 31575 14373 31609
rect 14239 31541 14289 31575
rect 14323 31541 14373 31575
rect 14239 31507 14373 31541
rect 14239 31473 14289 31507
rect 14323 31473 14373 31507
rect 14239 31439 14373 31473
rect 14239 31405 14289 31439
rect 14323 31405 14373 31439
rect 14239 31371 14373 31405
rect 14239 31337 14289 31371
rect 14323 31337 14373 31371
rect 14239 31303 14373 31337
rect 14239 31269 14289 31303
rect 14323 31269 14373 31303
rect 14239 31235 14373 31269
rect 14239 31201 14289 31235
rect 14323 31201 14373 31235
rect 14239 31167 14373 31201
rect 14239 31133 14289 31167
rect 14323 31133 14373 31167
rect 14239 31099 14373 31133
rect 14239 31065 14289 31099
rect 14323 31065 14373 31099
rect 14239 31031 14373 31065
rect 14239 30997 14289 31031
rect 14323 30997 14373 31031
rect 14239 30963 14373 30997
rect 14239 30929 14289 30963
rect 14323 30929 14373 30963
rect 14239 30895 14373 30929
rect 14239 30861 14289 30895
rect 14323 30861 14373 30895
rect 14239 30827 14373 30861
rect 14239 30793 14289 30827
rect 14323 30793 14373 30827
rect 14239 30759 14373 30793
rect 14239 30725 14289 30759
rect 14323 30725 14373 30759
rect 14239 30691 14373 30725
rect 14239 30657 14289 30691
rect 14323 30657 14373 30691
rect 14239 30623 14373 30657
rect 14239 30589 14289 30623
rect 14323 30589 14373 30623
rect 14239 30555 14373 30589
rect 14239 30521 14289 30555
rect 14323 30521 14373 30555
rect 14239 30487 14373 30521
rect 14239 30453 14289 30487
rect 14323 30453 14373 30487
rect 14239 30419 14373 30453
rect 14239 30385 14289 30419
rect 14323 30385 14373 30419
rect 14239 30351 14373 30385
rect 14239 30317 14289 30351
rect 14323 30317 14373 30351
rect 14239 30283 14373 30317
rect 14239 30249 14289 30283
rect 14323 30249 14373 30283
rect 14239 30215 14373 30249
rect 14239 30181 14289 30215
rect 14323 30181 14373 30215
rect 14239 30147 14373 30181
rect 14239 30113 14289 30147
rect 14323 30113 14373 30147
rect 14239 30079 14373 30113
rect 14239 30045 14289 30079
rect 14323 30045 14373 30079
rect 14239 30011 14373 30045
rect 14239 29977 14289 30011
rect 14323 29977 14373 30011
rect 14239 29943 14373 29977
rect 14239 29909 14289 29943
rect 14323 29909 14373 29943
rect 14239 29875 14373 29909
rect 14239 29841 14289 29875
rect 14323 29841 14373 29875
rect 14239 29807 14373 29841
rect 14239 29773 14289 29807
rect 14323 29773 14373 29807
rect 14239 29739 14373 29773
rect 14239 29705 14289 29739
rect 14323 29705 14373 29739
rect 14239 29671 14373 29705
rect 14239 29637 14289 29671
rect 14323 29637 14373 29671
rect 14239 29603 14373 29637
rect 14239 29569 14289 29603
rect 14323 29569 14373 29603
rect 14239 29535 14373 29569
rect 14239 29501 14289 29535
rect 14323 29501 14373 29535
rect 14239 29467 14373 29501
rect 14239 29433 14289 29467
rect 14323 29433 14373 29467
rect 14239 29399 14373 29433
rect 14239 29365 14289 29399
rect 14323 29365 14373 29399
rect 14239 29331 14373 29365
rect 14239 29297 14289 29331
rect 14323 29297 14373 29331
rect 14239 29263 14373 29297
rect 14239 29229 14289 29263
rect 14323 29229 14373 29263
rect 14239 29195 14373 29229
rect 14239 29161 14289 29195
rect 14323 29161 14373 29195
rect 14239 29127 14373 29161
rect 14239 29093 14289 29127
rect 14323 29093 14373 29127
rect 14239 29059 14373 29093
rect 14239 29025 14289 29059
rect 14323 29025 14373 29059
rect 14239 28991 14373 29025
rect 14239 28957 14289 28991
rect 14323 28957 14373 28991
rect 14239 28923 14373 28957
rect 14239 28889 14289 28923
rect 14323 28889 14373 28923
rect 14239 28855 14373 28889
rect 14239 28821 14289 28855
rect 14323 28821 14373 28855
rect 14239 28787 14373 28821
rect 14239 28753 14289 28787
rect 14323 28753 14373 28787
rect 14239 28719 14373 28753
rect 14239 28685 14289 28719
rect 14323 28685 14373 28719
rect 14239 28651 14373 28685
rect 14239 28617 14289 28651
rect 14323 28617 14373 28651
rect 14239 28583 14373 28617
rect 14239 28549 14289 28583
rect 14323 28549 14373 28583
rect 14239 28515 14373 28549
rect 14239 28481 14289 28515
rect 14323 28481 14373 28515
rect 14239 28447 14373 28481
rect 14239 28413 14289 28447
rect 14323 28413 14373 28447
rect 14239 28379 14373 28413
rect 14239 28345 14289 28379
rect 14323 28345 14373 28379
rect 14239 28311 14373 28345
rect 14239 28277 14289 28311
rect 14323 28277 14373 28311
rect 14239 28243 14373 28277
rect 14239 28209 14289 28243
rect 14323 28209 14373 28243
rect 14239 28175 14373 28209
rect 14239 28141 14289 28175
rect 14323 28141 14373 28175
rect 14239 28107 14373 28141
rect 14239 28073 14289 28107
rect 14323 28073 14373 28107
rect 14239 28039 14373 28073
rect 14239 28005 14289 28039
rect 14323 28005 14373 28039
rect 14239 27971 14373 28005
rect 14239 27937 14289 27971
rect 14323 27937 14373 27971
rect 14239 27903 14373 27937
rect 14239 27869 14289 27903
rect 14323 27869 14373 27903
rect 14239 27835 14373 27869
rect 14239 27801 14289 27835
rect 14323 27801 14373 27835
rect 14239 27767 14373 27801
rect 14239 27733 14289 27767
rect 14323 27733 14373 27767
rect 14239 27699 14373 27733
rect 14239 27665 14289 27699
rect 14323 27665 14373 27699
rect 14239 27631 14373 27665
rect 14239 27597 14289 27631
rect 14323 27597 14373 27631
rect 14239 27563 14373 27597
rect 14239 27529 14289 27563
rect 14323 27529 14373 27563
rect 14239 27495 14373 27529
rect 14239 27461 14289 27495
rect 14323 27461 14373 27495
rect 14239 27427 14373 27461
rect 14239 27393 14289 27427
rect 14323 27393 14373 27427
rect 14239 27359 14373 27393
rect 14239 27325 14289 27359
rect 14323 27325 14373 27359
rect 14239 27291 14373 27325
rect 14239 27257 14289 27291
rect 14323 27257 14373 27291
rect 14239 27223 14373 27257
rect 14239 27189 14289 27223
rect 14323 27189 14373 27223
rect 14239 27155 14373 27189
rect 14239 27121 14289 27155
rect 14323 27121 14373 27155
rect 14239 27087 14373 27121
rect 14239 27053 14289 27087
rect 14323 27053 14373 27087
rect 14239 27019 14373 27053
rect 14239 26985 14289 27019
rect 14323 26985 14373 27019
rect 14239 26951 14373 26985
rect 14239 26917 14289 26951
rect 14323 26917 14373 26951
rect 14239 26883 14373 26917
rect 14239 26849 14289 26883
rect 14323 26849 14373 26883
rect 14239 26815 14373 26849
rect 14239 26781 14289 26815
rect 14323 26781 14373 26815
rect 14239 26747 14373 26781
rect 14239 26713 14289 26747
rect 14323 26713 14373 26747
rect 14239 26679 14373 26713
rect 14239 26645 14289 26679
rect 14323 26645 14373 26679
rect 14239 26611 14373 26645
rect 14239 26577 14289 26611
rect 14323 26577 14373 26611
rect 14239 26543 14373 26577
rect 14239 26509 14289 26543
rect 14323 26509 14373 26543
rect 14239 26475 14373 26509
rect 14239 26441 14289 26475
rect 14323 26441 14373 26475
rect 14239 26407 14373 26441
rect 14239 26373 14289 26407
rect 14323 26373 14373 26407
rect 14239 26339 14373 26373
rect 14239 26305 14289 26339
rect 14323 26305 14373 26339
rect 14239 26271 14373 26305
rect 14239 26237 14289 26271
rect 14323 26237 14373 26271
rect 14239 26203 14373 26237
rect 14239 26169 14289 26203
rect 14323 26169 14373 26203
rect 14239 26135 14373 26169
rect 14239 26101 14289 26135
rect 14323 26101 14373 26135
rect 14239 26067 14373 26101
rect 14239 26033 14289 26067
rect 14323 26033 14373 26067
rect 14239 25999 14373 26033
rect 14239 25965 14289 25999
rect 14323 25965 14373 25999
rect 14239 25931 14373 25965
rect 14239 25897 14289 25931
rect 14323 25897 14373 25931
rect 14239 25863 14373 25897
rect 14239 25829 14289 25863
rect 14323 25829 14373 25863
rect 14239 25795 14373 25829
rect 14239 25761 14289 25795
rect 14323 25761 14373 25795
rect 14239 25727 14373 25761
rect 14239 25693 14289 25727
rect 14323 25693 14373 25727
rect 14239 25659 14373 25693
rect 14239 25625 14289 25659
rect 14323 25625 14373 25659
rect 14239 25591 14373 25625
rect 14239 25557 14289 25591
rect 14323 25557 14373 25591
rect 14239 25523 14373 25557
rect 14239 25489 14289 25523
rect 14323 25489 14373 25523
rect 14239 25455 14373 25489
rect 14239 25421 14289 25455
rect 14323 25421 14373 25455
rect 14239 25387 14373 25421
rect 14239 25353 14289 25387
rect 14323 25353 14373 25387
rect 14239 25319 14373 25353
rect 14239 25285 14289 25319
rect 14323 25285 14373 25319
rect 14239 25251 14373 25285
rect 14239 25217 14289 25251
rect 14323 25217 14373 25251
rect 14239 25183 14373 25217
rect 14239 25149 14289 25183
rect 14323 25149 14373 25183
rect 14239 25115 14373 25149
rect 14239 25081 14289 25115
rect 14323 25081 14373 25115
rect 14239 25047 14373 25081
rect 14239 25013 14289 25047
rect 14323 25013 14373 25047
rect 14239 24979 14373 25013
rect 14239 24945 14289 24979
rect 14323 24945 14373 24979
rect 14239 24911 14373 24945
rect 14239 24877 14289 24911
rect 14323 24877 14373 24911
rect 14239 24843 14373 24877
rect 14239 24809 14289 24843
rect 14323 24809 14373 24843
rect 14239 24775 14373 24809
rect 14239 24741 14289 24775
rect 14323 24741 14373 24775
rect 14239 24707 14373 24741
rect 14239 24673 14289 24707
rect 14323 24673 14373 24707
rect 14239 24639 14373 24673
rect 14239 24605 14289 24639
rect 14323 24605 14373 24639
rect 14239 24571 14373 24605
rect 14239 24537 14289 24571
rect 14323 24537 14373 24571
rect 14239 24503 14373 24537
rect 14239 24469 14289 24503
rect 14323 24469 14373 24503
rect 14239 24435 14373 24469
rect 14239 24401 14289 24435
rect 14323 24401 14373 24435
rect 14239 24367 14373 24401
rect 14239 24333 14289 24367
rect 14323 24333 14373 24367
rect 14239 24299 14373 24333
rect 14239 24265 14289 24299
rect 14323 24265 14373 24299
rect 14239 24231 14373 24265
rect 14239 24197 14289 24231
rect 14323 24197 14373 24231
rect 14239 24163 14373 24197
rect 14239 24129 14289 24163
rect 14323 24129 14373 24163
rect 14239 24095 14373 24129
rect 14239 24061 14289 24095
rect 14323 24061 14373 24095
rect 14239 24027 14373 24061
rect 14239 23993 14289 24027
rect 14323 23993 14373 24027
rect 14239 23959 14373 23993
rect 14239 23925 14289 23959
rect 14323 23925 14373 23959
rect 14239 23891 14373 23925
rect 14239 23857 14289 23891
rect 14323 23857 14373 23891
rect 14239 23823 14373 23857
rect 14239 23789 14289 23823
rect 14323 23789 14373 23823
rect 14239 23755 14373 23789
rect 14239 23721 14289 23755
rect 14323 23721 14373 23755
rect 14239 23687 14373 23721
rect 14239 23653 14289 23687
rect 14323 23653 14373 23687
rect 14239 23619 14373 23653
rect 14239 23585 14289 23619
rect 14323 23585 14373 23619
rect 14239 23551 14373 23585
rect 14239 23517 14289 23551
rect 14323 23517 14373 23551
rect 14239 23483 14373 23517
rect 14239 23449 14289 23483
rect 14323 23449 14373 23483
rect 14239 23415 14373 23449
rect 14239 23381 14289 23415
rect 14323 23381 14373 23415
rect 14239 23347 14373 23381
rect 14239 23313 14289 23347
rect 14323 23313 14373 23347
rect 14239 23279 14373 23313
rect 14239 23245 14289 23279
rect 14323 23245 14373 23279
rect 14239 23211 14373 23245
rect 14239 23177 14289 23211
rect 14323 23177 14373 23211
rect 14239 23143 14373 23177
rect 14239 23109 14289 23143
rect 14323 23109 14373 23143
rect 14239 23075 14373 23109
rect 14239 23041 14289 23075
rect 14323 23041 14373 23075
rect 14239 23007 14373 23041
rect 14239 22973 14289 23007
rect 14323 22973 14373 23007
rect 14239 22939 14373 22973
rect 14239 22905 14289 22939
rect 14323 22905 14373 22939
rect 14239 22871 14373 22905
rect 14239 22837 14289 22871
rect 14323 22837 14373 22871
rect 14239 22803 14373 22837
rect 14239 22769 14289 22803
rect 14323 22769 14373 22803
rect 14239 22735 14373 22769
rect 14239 22701 14289 22735
rect 14323 22701 14373 22735
rect 14239 22667 14373 22701
rect 14239 22633 14289 22667
rect 14323 22633 14373 22667
rect 14239 22599 14373 22633
rect 14239 22565 14289 22599
rect 14323 22565 14373 22599
rect 14239 22531 14373 22565
rect 14239 22497 14289 22531
rect 14323 22497 14373 22531
rect 14239 22463 14373 22497
rect 14239 22429 14289 22463
rect 14323 22429 14373 22463
rect 14239 22395 14373 22429
rect 14239 22361 14289 22395
rect 14323 22361 14373 22395
rect 14239 22327 14373 22361
rect 14239 22293 14289 22327
rect 14323 22293 14373 22327
rect 14239 22259 14373 22293
rect 14239 22225 14289 22259
rect 14323 22225 14373 22259
rect 14239 22191 14373 22225
rect 14239 22157 14289 22191
rect 14323 22157 14373 22191
rect 14239 22123 14373 22157
rect 14239 22089 14289 22123
rect 14323 22089 14373 22123
rect 14239 22055 14373 22089
rect 14239 22021 14289 22055
rect 14323 22021 14373 22055
rect 14239 21987 14373 22021
rect 14239 21953 14289 21987
rect 14323 21953 14373 21987
rect 14239 21919 14373 21953
rect 14239 21885 14289 21919
rect 14323 21885 14373 21919
rect 14239 21851 14373 21885
rect 14239 21817 14289 21851
rect 14323 21817 14373 21851
rect 14239 21783 14373 21817
rect 14239 21749 14289 21783
rect 14323 21749 14373 21783
rect 14239 21715 14373 21749
rect 14239 21681 14289 21715
rect 14323 21681 14373 21715
rect 14239 21647 14373 21681
rect 14239 21613 14289 21647
rect 14323 21613 14373 21647
rect 14239 21579 14373 21613
rect 14239 21545 14289 21579
rect 14323 21545 14373 21579
rect 14239 21511 14373 21545
rect 14239 21477 14289 21511
rect 14323 21477 14373 21511
rect 14239 21443 14373 21477
rect 14239 21409 14289 21443
rect 14323 21409 14373 21443
rect 14239 21375 14373 21409
rect 14239 21341 14289 21375
rect 14323 21341 14373 21375
rect 14239 21307 14373 21341
rect 14239 21273 14289 21307
rect 14323 21273 14373 21307
rect 14239 21239 14373 21273
rect 14239 21205 14289 21239
rect 14323 21205 14373 21239
rect 14239 21171 14373 21205
rect 14239 21137 14289 21171
rect 14323 21137 14373 21171
rect 14239 21103 14373 21137
rect 14239 21069 14289 21103
rect 14323 21069 14373 21103
rect 14239 21035 14373 21069
rect 14239 21001 14289 21035
rect 14323 21001 14373 21035
rect 14239 20967 14373 21001
rect 14239 20933 14289 20967
rect 14323 20933 14373 20967
rect 14239 20899 14373 20933
rect 14239 20865 14289 20899
rect 14323 20865 14373 20899
rect 14239 20831 14373 20865
rect 14239 20797 14289 20831
rect 14323 20797 14373 20831
rect 14239 20763 14373 20797
rect 14239 20729 14289 20763
rect 14323 20729 14373 20763
rect 14239 20695 14373 20729
rect 14239 20661 14289 20695
rect 14323 20661 14373 20695
rect 14239 20627 14373 20661
rect 14239 20593 14289 20627
rect 14323 20593 14373 20627
rect 14239 20559 14373 20593
rect 14239 20525 14289 20559
rect 14323 20525 14373 20559
rect 14239 20491 14373 20525
rect 14239 20457 14289 20491
rect 14323 20457 14373 20491
rect 14239 20423 14373 20457
rect 14239 20389 14289 20423
rect 14323 20389 14373 20423
rect 14239 20355 14373 20389
rect 14239 20321 14289 20355
rect 14323 20321 14373 20355
rect 14239 20287 14373 20321
rect 14239 20253 14289 20287
rect 14323 20253 14373 20287
rect 14239 20219 14373 20253
rect 14239 20185 14289 20219
rect 14323 20185 14373 20219
rect 14239 20151 14373 20185
rect 14239 20117 14289 20151
rect 14323 20117 14373 20151
rect 14239 20083 14373 20117
rect 14239 20049 14289 20083
rect 14323 20049 14373 20083
rect 14239 20015 14373 20049
rect 14239 19981 14289 20015
rect 14323 19981 14373 20015
rect 14239 19947 14373 19981
rect 14239 19913 14289 19947
rect 14323 19913 14373 19947
rect 14239 19879 14373 19913
rect 14239 19845 14289 19879
rect 14323 19845 14373 19879
rect 14239 19811 14373 19845
rect 14239 19777 14289 19811
rect 14323 19777 14373 19811
rect 14239 19743 14373 19777
rect 14239 19709 14289 19743
rect 14323 19709 14373 19743
rect 14239 19675 14373 19709
rect 14239 19641 14289 19675
rect 14323 19641 14373 19675
rect 14239 19607 14373 19641
rect 14239 19573 14289 19607
rect 14323 19573 14373 19607
rect 14239 19539 14373 19573
rect 14239 19505 14289 19539
rect 14323 19505 14373 19539
rect 14239 19471 14373 19505
rect 14239 19437 14289 19471
rect 14323 19437 14373 19471
rect 14239 19403 14373 19437
rect 14239 19369 14289 19403
rect 14323 19369 14373 19403
rect 14239 19335 14373 19369
rect 14239 19301 14289 19335
rect 14323 19301 14373 19335
rect 14239 19267 14373 19301
rect 14239 19233 14289 19267
rect 14323 19233 14373 19267
rect 14239 19199 14373 19233
rect 14239 19165 14289 19199
rect 14323 19165 14373 19199
rect 14239 19131 14373 19165
rect 14239 19097 14289 19131
rect 14323 19097 14373 19131
rect 14239 19063 14373 19097
rect 14239 19029 14289 19063
rect 14323 19029 14373 19063
rect 14239 18995 14373 19029
rect 14239 18961 14289 18995
rect 14323 18961 14373 18995
rect 14239 18927 14373 18961
rect 14239 18893 14289 18927
rect 14323 18893 14373 18927
rect 14239 18859 14373 18893
rect 14239 18825 14289 18859
rect 14323 18825 14373 18859
rect 14239 18791 14373 18825
rect 14239 18757 14289 18791
rect 14323 18757 14373 18791
rect 14239 18723 14373 18757
rect 14239 18689 14289 18723
rect 14323 18689 14373 18723
rect 14239 18655 14373 18689
rect 14239 18621 14289 18655
rect 14323 18621 14373 18655
rect 14239 18587 14373 18621
rect 14239 18553 14289 18587
rect 14323 18553 14373 18587
rect 14239 18519 14373 18553
rect 14239 18485 14289 18519
rect 14323 18485 14373 18519
rect 14239 18451 14373 18485
rect 14239 18417 14289 18451
rect 14323 18417 14373 18451
rect 14239 18383 14373 18417
rect 14239 18349 14289 18383
rect 14323 18349 14373 18383
rect 14239 18315 14373 18349
rect 14239 18281 14289 18315
rect 14323 18281 14373 18315
rect 14239 18247 14373 18281
rect 14239 18213 14289 18247
rect 14323 18213 14373 18247
rect 14239 18179 14373 18213
rect 14239 18145 14289 18179
rect 14323 18145 14373 18179
rect 14239 18111 14373 18145
rect 14239 18077 14289 18111
rect 14323 18077 14373 18111
rect 14239 18043 14373 18077
rect 14239 18009 14289 18043
rect 14323 18009 14373 18043
rect 14239 17975 14373 18009
rect 14239 17941 14289 17975
rect 14323 17941 14373 17975
rect 14239 17907 14373 17941
rect 14239 17873 14289 17907
rect 14323 17873 14373 17907
rect 14239 17839 14373 17873
rect 14239 17805 14289 17839
rect 14323 17805 14373 17839
rect 14239 17771 14373 17805
rect 14239 17737 14289 17771
rect 14323 17737 14373 17771
rect 14239 17703 14373 17737
rect 14239 17669 14289 17703
rect 14323 17669 14373 17703
rect 14239 17635 14373 17669
rect 14239 17601 14289 17635
rect 14323 17601 14373 17635
rect 14239 17567 14373 17601
rect 14239 17533 14289 17567
rect 14323 17533 14373 17567
rect 14239 17499 14373 17533
rect 14239 17465 14289 17499
rect 14323 17465 14373 17499
rect 14239 17431 14373 17465
rect 14239 17397 14289 17431
rect 14323 17397 14373 17431
rect 14239 17363 14373 17397
rect 14239 17329 14289 17363
rect 14323 17329 14373 17363
rect 14239 17295 14373 17329
rect 14239 17261 14289 17295
rect 14323 17261 14373 17295
rect 14239 17227 14373 17261
rect 14239 17193 14289 17227
rect 14323 17193 14373 17227
rect 14239 17159 14373 17193
rect 14239 17125 14289 17159
rect 14323 17125 14373 17159
rect 14239 17091 14373 17125
rect 14239 17057 14289 17091
rect 14323 17057 14373 17091
rect 14239 17023 14373 17057
rect 14239 16989 14289 17023
rect 14323 16989 14373 17023
rect 14239 16955 14373 16989
rect 14239 16921 14289 16955
rect 14323 16921 14373 16955
rect 14239 16887 14373 16921
rect 14239 16853 14289 16887
rect 14323 16853 14373 16887
rect 14239 16819 14373 16853
rect 14239 16785 14289 16819
rect 14323 16785 14373 16819
rect 14239 16751 14373 16785
rect 14239 16717 14289 16751
rect 14323 16717 14373 16751
rect 14239 16683 14373 16717
rect 14239 16649 14289 16683
rect 14323 16649 14373 16683
rect 14239 16615 14373 16649
rect 14239 16581 14289 16615
rect 14323 16581 14373 16615
rect 14239 16547 14373 16581
rect 14239 16513 14289 16547
rect 14323 16513 14373 16547
rect 14239 16479 14373 16513
rect 14239 16445 14289 16479
rect 14323 16445 14373 16479
rect 14239 16411 14373 16445
rect 14239 16377 14289 16411
rect 14323 16377 14373 16411
rect 14239 16343 14373 16377
rect 14239 16309 14289 16343
rect 14323 16309 14373 16343
rect 14239 16275 14373 16309
rect 14239 16241 14289 16275
rect 14323 16241 14373 16275
rect 14239 16207 14373 16241
rect 14239 16173 14289 16207
rect 14323 16173 14373 16207
rect 14239 16139 14373 16173
rect 14239 16105 14289 16139
rect 14323 16105 14373 16139
rect 14239 16071 14373 16105
rect 14239 16037 14289 16071
rect 14323 16037 14373 16071
rect 14239 16003 14373 16037
rect 14239 15969 14289 16003
rect 14323 15969 14373 16003
rect 14239 15935 14373 15969
rect 14239 15901 14289 15935
rect 14323 15901 14373 15935
rect 14239 15867 14373 15901
rect 14239 15833 14289 15867
rect 14323 15833 14373 15867
rect 14239 15799 14373 15833
rect 14239 15765 14289 15799
rect 14323 15765 14373 15799
rect 14239 15731 14373 15765
rect 14239 15697 14289 15731
rect 14323 15697 14373 15731
rect 14239 15663 14373 15697
rect 14239 15629 14289 15663
rect 14323 15629 14373 15663
rect 14239 15595 14373 15629
rect 14239 15561 14289 15595
rect 14323 15561 14373 15595
rect 14239 15527 14373 15561
rect 14239 15493 14289 15527
rect 14323 15493 14373 15527
rect 14239 15459 14373 15493
rect 14239 15425 14289 15459
rect 14323 15425 14373 15459
rect 14239 15391 14373 15425
rect 14239 15357 14289 15391
rect 14323 15357 14373 15391
rect 14239 15323 14373 15357
rect 14239 15289 14289 15323
rect 14323 15289 14373 15323
rect 14239 15255 14373 15289
rect 14239 15221 14289 15255
rect 14323 15221 14373 15255
rect 575 15153 624 15187
rect 658 15153 707 15187
rect 575 15119 707 15153
rect 575 15085 624 15119
rect 658 15085 707 15119
rect 575 15051 707 15085
rect 575 15017 624 15051
rect 658 15017 707 15051
rect 575 14983 707 15017
rect 575 14949 624 14983
rect 658 14949 707 14983
rect 575 14915 707 14949
rect 575 14881 624 14915
rect 658 14881 707 14915
rect 575 14838 707 14881
rect 14239 15187 14373 15221
rect 14239 15153 14289 15187
rect 14323 15153 14373 15187
rect 14239 15119 14373 15153
rect 14239 15085 14289 15119
rect 14323 15085 14373 15119
rect 14239 15051 14373 15085
rect 14239 15017 14289 15051
rect 14323 15017 14373 15051
rect 14239 14983 14373 15017
rect 14239 14949 14289 14983
rect 14323 14949 14373 14983
rect 14239 14915 14373 14949
rect 14239 14881 14289 14915
rect 14323 14881 14373 14915
rect 14239 14838 14373 14881
rect 575 14788 14373 14838
rect 575 14754 758 14788
rect 792 14754 826 14788
rect 860 14754 894 14788
rect 928 14754 962 14788
rect 996 14754 1030 14788
rect 1064 14754 1098 14788
rect 1132 14754 1166 14788
rect 1200 14754 1234 14788
rect 1268 14754 1302 14788
rect 1336 14754 1370 14788
rect 1404 14754 1438 14788
rect 1472 14754 1506 14788
rect 1540 14754 1574 14788
rect 1608 14754 1642 14788
rect 1676 14754 1710 14788
rect 1744 14754 1778 14788
rect 1812 14754 1846 14788
rect 1880 14754 1914 14788
rect 1948 14754 1982 14788
rect 2016 14754 2050 14788
rect 2084 14754 2118 14788
rect 2152 14754 2186 14788
rect 2220 14754 2254 14788
rect 2288 14754 2322 14788
rect 2356 14754 2390 14788
rect 2424 14754 2458 14788
rect 2492 14754 2526 14788
rect 2560 14754 2594 14788
rect 2628 14754 2662 14788
rect 2696 14754 2730 14788
rect 2764 14754 2798 14788
rect 2832 14754 2866 14788
rect 2900 14754 2934 14788
rect 2968 14754 3002 14788
rect 3036 14754 3070 14788
rect 3104 14754 3138 14788
rect 3172 14754 3206 14788
rect 3240 14754 3274 14788
rect 3308 14754 3342 14788
rect 3376 14754 3410 14788
rect 3444 14754 3478 14788
rect 3512 14754 3546 14788
rect 3580 14754 3614 14788
rect 3648 14754 3682 14788
rect 3716 14754 3750 14788
rect 3784 14754 3818 14788
rect 3852 14754 3886 14788
rect 3920 14754 3954 14788
rect 3988 14754 4022 14788
rect 4056 14754 4090 14788
rect 4124 14754 4158 14788
rect 4192 14754 4226 14788
rect 4260 14754 4294 14788
rect 4328 14754 4362 14788
rect 4396 14754 4430 14788
rect 4464 14754 4498 14788
rect 4532 14754 4566 14788
rect 4600 14754 4634 14788
rect 4668 14754 4702 14788
rect 4736 14754 4770 14788
rect 4804 14754 4838 14788
rect 4872 14754 4906 14788
rect 4940 14754 4974 14788
rect 5008 14754 5042 14788
rect 5076 14754 5110 14788
rect 5144 14754 5178 14788
rect 5212 14754 5246 14788
rect 5280 14754 5314 14788
rect 5348 14754 5382 14788
rect 5416 14754 5450 14788
rect 5484 14754 5518 14788
rect 5552 14754 5586 14788
rect 5620 14754 5654 14788
rect 5688 14754 5722 14788
rect 5756 14754 5790 14788
rect 5824 14754 5858 14788
rect 5892 14754 5926 14788
rect 5960 14754 5994 14788
rect 6028 14754 6062 14788
rect 6096 14754 6130 14788
rect 6164 14754 6198 14788
rect 6232 14754 6266 14788
rect 6300 14754 6334 14788
rect 6368 14754 6402 14788
rect 6436 14754 6470 14788
rect 6504 14754 6538 14788
rect 6572 14754 6606 14788
rect 6640 14754 6674 14788
rect 6708 14754 6742 14788
rect 6776 14754 6810 14788
rect 6844 14754 6878 14788
rect 6912 14754 6946 14788
rect 6980 14754 7014 14788
rect 7048 14754 7082 14788
rect 7116 14754 7150 14788
rect 7184 14754 7218 14788
rect 7252 14754 7286 14788
rect 7320 14754 7354 14788
rect 7388 14754 7422 14788
rect 7456 14754 7490 14788
rect 7524 14754 7558 14788
rect 7592 14754 7626 14788
rect 7660 14754 7694 14788
rect 7728 14754 7762 14788
rect 7796 14754 7830 14788
rect 7864 14754 7898 14788
rect 7932 14754 7966 14788
rect 8000 14754 8034 14788
rect 8068 14754 8102 14788
rect 8136 14754 8170 14788
rect 8204 14754 8238 14788
rect 8272 14754 8306 14788
rect 8340 14754 8374 14788
rect 8408 14754 8442 14788
rect 8476 14754 8510 14788
rect 8544 14754 8578 14788
rect 8612 14754 8646 14788
rect 8680 14754 8714 14788
rect 8748 14754 8782 14788
rect 8816 14754 8850 14788
rect 8884 14754 8918 14788
rect 8952 14754 8986 14788
rect 9020 14754 9054 14788
rect 9088 14754 9122 14788
rect 9156 14754 9190 14788
rect 9224 14754 9258 14788
rect 9292 14754 9326 14788
rect 9360 14754 9394 14788
rect 9428 14754 9462 14788
rect 9496 14754 9530 14788
rect 9564 14754 9598 14788
rect 9632 14754 9666 14788
rect 9700 14754 9734 14788
rect 9768 14754 9802 14788
rect 9836 14754 9870 14788
rect 9904 14754 9938 14788
rect 9972 14754 10006 14788
rect 10040 14754 10074 14788
rect 10108 14754 10142 14788
rect 10176 14754 10210 14788
rect 10244 14754 10278 14788
rect 10312 14754 10346 14788
rect 10380 14754 10414 14788
rect 10448 14754 10482 14788
rect 10516 14754 10550 14788
rect 10584 14754 10618 14788
rect 10652 14754 10686 14788
rect 10720 14754 10754 14788
rect 10788 14754 10822 14788
rect 10856 14754 10890 14788
rect 10924 14754 10958 14788
rect 10992 14754 11026 14788
rect 11060 14754 11094 14788
rect 11128 14754 11162 14788
rect 11196 14754 11230 14788
rect 11264 14754 11298 14788
rect 11332 14754 11366 14788
rect 11400 14754 11434 14788
rect 11468 14754 11502 14788
rect 11536 14754 11570 14788
rect 11604 14754 11638 14788
rect 11672 14754 11706 14788
rect 11740 14754 11774 14788
rect 11808 14754 11842 14788
rect 11876 14754 11910 14788
rect 11944 14754 11978 14788
rect 12012 14754 12046 14788
rect 12080 14754 12114 14788
rect 12148 14754 12182 14788
rect 12216 14754 12250 14788
rect 12284 14754 12318 14788
rect 12352 14754 12386 14788
rect 12420 14754 12454 14788
rect 12488 14754 12522 14788
rect 12556 14754 12590 14788
rect 12624 14754 12658 14788
rect 12692 14754 12726 14788
rect 12760 14754 12794 14788
rect 12828 14754 12862 14788
rect 12896 14754 12930 14788
rect 12964 14754 12998 14788
rect 13032 14754 13066 14788
rect 13100 14754 13134 14788
rect 13168 14754 13202 14788
rect 13236 14754 13270 14788
rect 13304 14754 13338 14788
rect 13372 14754 13406 14788
rect 13440 14754 13474 14788
rect 13508 14754 13542 14788
rect 13576 14754 13610 14788
rect 13644 14754 13678 14788
rect 13712 14754 13746 14788
rect 13780 14754 13814 14788
rect 13848 14754 13882 14788
rect 13916 14754 13950 14788
rect 13984 14754 14018 14788
rect 14052 14754 14086 14788
rect 14120 14754 14154 14788
rect 14188 14754 14373 14788
rect 575 14704 14373 14754
<< mvpsubdiffcont >>
rect 447 36476 481 36510
rect 515 36476 549 36510
rect 583 36476 617 36510
rect 651 36476 685 36510
rect 719 36476 753 36510
rect 787 36476 821 36510
rect 855 36476 889 36510
rect 923 36476 957 36510
rect 991 36476 1025 36510
rect 1059 36476 1093 36510
rect 1127 36476 1161 36510
rect 1195 36476 1229 36510
rect 1263 36476 1297 36510
rect 1331 36476 1365 36510
rect 1399 36476 1433 36510
rect 1467 36476 1501 36510
rect 1535 36476 1569 36510
rect 1603 36476 1637 36510
rect 1671 36476 1705 36510
rect 1739 36476 1773 36510
rect 1807 36476 1841 36510
rect 1875 36476 1909 36510
rect 1943 36476 1977 36510
rect 2011 36476 2045 36510
rect 2079 36476 2113 36510
rect 2147 36476 2181 36510
rect 2215 36476 2249 36510
rect 2283 36476 2317 36510
rect 2351 36476 2385 36510
rect 2419 36476 2453 36510
rect 2487 36476 2521 36510
rect 2555 36476 2589 36510
rect 2623 36476 2657 36510
rect 2691 36476 2725 36510
rect 2759 36476 2793 36510
rect 2827 36476 2861 36510
rect 2895 36476 2929 36510
rect 2963 36476 2997 36510
rect 3031 36476 3065 36510
rect 3099 36476 3133 36510
rect 3167 36476 3201 36510
rect 3235 36476 3269 36510
rect 3303 36476 3337 36510
rect 3371 36476 3405 36510
rect 3439 36476 3473 36510
rect 3507 36476 3541 36510
rect 3575 36476 3609 36510
rect 3643 36476 3677 36510
rect 3711 36476 3745 36510
rect 3779 36476 3813 36510
rect 3847 36476 3881 36510
rect 3915 36476 3949 36510
rect 3983 36476 4017 36510
rect 4051 36476 4085 36510
rect 4119 36476 4153 36510
rect 4187 36476 4221 36510
rect 4255 36476 4289 36510
rect 4323 36476 4357 36510
rect 4391 36476 4425 36510
rect 4459 36476 4493 36510
rect 4527 36476 4561 36510
rect 4595 36476 4629 36510
rect 4663 36476 4697 36510
rect 4731 36476 4765 36510
rect 4799 36476 4833 36510
rect 4867 36476 4901 36510
rect 4935 36476 4969 36510
rect 5003 36476 5037 36510
rect 5071 36476 5105 36510
rect 5139 36476 5173 36510
rect 5207 36476 5241 36510
rect 5275 36476 5309 36510
rect 5343 36476 5377 36510
rect 5411 36476 5445 36510
rect 5479 36476 5513 36510
rect 5547 36476 5581 36510
rect 5615 36476 5649 36510
rect 5683 36476 5717 36510
rect 5751 36476 5785 36510
rect 5819 36476 5853 36510
rect 5887 36476 5921 36510
rect 5955 36476 5989 36510
rect 6023 36476 6057 36510
rect 6091 36476 6125 36510
rect 6159 36476 6193 36510
rect 6227 36476 6261 36510
rect 6295 36476 6329 36510
rect 6363 36476 6397 36510
rect 6431 36476 6465 36510
rect 6499 36476 6533 36510
rect 6567 36476 6601 36510
rect 6635 36476 6669 36510
rect 6703 36476 6737 36510
rect 6771 36476 6805 36510
rect 6839 36476 6873 36510
rect 6907 36476 6941 36510
rect 6975 36476 7009 36510
rect 7043 36476 7077 36510
rect 7111 36476 7145 36510
rect 7179 36476 7213 36510
rect 7247 36476 7281 36510
rect 7315 36476 7349 36510
rect 7383 36476 7417 36510
rect 7451 36476 7485 36510
rect 7519 36476 7553 36510
rect 7587 36476 7621 36510
rect 7655 36476 7689 36510
rect 7723 36476 7757 36510
rect 7791 36476 7825 36510
rect 7859 36476 7893 36510
rect 7927 36476 7961 36510
rect 7995 36476 8029 36510
rect 8063 36476 8097 36510
rect 8131 36476 8165 36510
rect 8199 36476 8233 36510
rect 8267 36476 8301 36510
rect 8335 36476 8369 36510
rect 8403 36476 8437 36510
rect 8471 36476 8505 36510
rect 8539 36476 8573 36510
rect 8607 36476 8641 36510
rect 8675 36476 8709 36510
rect 8743 36476 8777 36510
rect 8811 36476 8845 36510
rect 8879 36476 8913 36510
rect 8947 36476 8981 36510
rect 9015 36476 9049 36510
rect 9083 36476 9117 36510
rect 9151 36476 9185 36510
rect 9219 36476 9253 36510
rect 9287 36476 9321 36510
rect 9355 36476 9389 36510
rect 9423 36476 9457 36510
rect 9491 36476 9525 36510
rect 9559 36476 9593 36510
rect 9627 36476 9661 36510
rect 9695 36476 9729 36510
rect 9763 36476 9797 36510
rect 9831 36476 9865 36510
rect 9899 36476 9933 36510
rect 9967 36476 10001 36510
rect 10035 36476 10069 36510
rect 10103 36476 10137 36510
rect 10171 36476 10205 36510
rect 10239 36476 10273 36510
rect 10307 36476 10341 36510
rect 10375 36476 10409 36510
rect 10443 36476 10477 36510
rect 10511 36476 10545 36510
rect 10579 36476 10613 36510
rect 10647 36476 10681 36510
rect 10715 36476 10749 36510
rect 10783 36476 10817 36510
rect 10851 36476 10885 36510
rect 10919 36476 10953 36510
rect 10987 36476 11021 36510
rect 11055 36476 11089 36510
rect 11123 36476 11157 36510
rect 11191 36476 11225 36510
rect 11259 36476 11293 36510
rect 11327 36476 11361 36510
rect 11395 36476 11429 36510
rect 11463 36476 11497 36510
rect 11531 36476 11565 36510
rect 11599 36476 11633 36510
rect 11667 36476 11701 36510
rect 11735 36476 11769 36510
rect 11803 36476 11837 36510
rect 11871 36476 11905 36510
rect 11939 36476 11973 36510
rect 12007 36476 12041 36510
rect 12075 36476 12109 36510
rect 12143 36476 12177 36510
rect 12211 36476 12245 36510
rect 12279 36476 12313 36510
rect 12347 36476 12381 36510
rect 12415 36476 12449 36510
rect 12483 36476 12517 36510
rect 12551 36476 12585 36510
rect 12619 36476 12653 36510
rect 12687 36476 12721 36510
rect 12755 36476 12789 36510
rect 12823 36476 12857 36510
rect 12891 36476 12925 36510
rect 12959 36476 12993 36510
rect 13027 36476 13061 36510
rect 13095 36476 13129 36510
rect 13163 36476 13197 36510
rect 13231 36476 13265 36510
rect 13299 36476 13333 36510
rect 13367 36476 13401 36510
rect 13435 36476 13469 36510
rect 13503 36476 13537 36510
rect 13571 36476 13605 36510
rect 13639 36476 13673 36510
rect 13707 36476 13741 36510
rect 13775 36476 13809 36510
rect 13843 36476 13877 36510
rect 13911 36476 13945 36510
rect 13979 36476 14013 36510
rect 14047 36476 14081 36510
rect 14115 36476 14149 36510
rect 14183 36476 14217 36510
rect 14251 36476 14285 36510
rect 14319 36476 14353 36510
rect 14387 36476 14421 36510
rect 14455 36476 14489 36510
rect 304 36335 338 36369
rect 304 36267 338 36301
rect 14599 36341 14633 36375
rect 14599 36273 14633 36307
rect 304 36199 338 36233
rect 304 36131 338 36165
rect 304 36063 338 36097
rect 304 35995 338 36029
rect 304 35927 338 35961
rect 304 35859 338 35893
rect 304 35791 338 35825
rect 304 35723 338 35757
rect 304 35655 338 35689
rect 304 35587 338 35621
rect 304 35519 338 35553
rect 304 35451 338 35485
rect 304 35383 338 35417
rect 304 35315 338 35349
rect 304 35247 338 35281
rect 304 35179 338 35213
rect 304 35111 338 35145
rect 304 35043 338 35077
rect 304 34975 338 35009
rect 304 34907 338 34941
rect 304 34839 338 34873
rect 304 34771 338 34805
rect 304 34703 338 34737
rect 304 34635 338 34669
rect 304 34567 338 34601
rect 304 34499 338 34533
rect 304 34431 338 34465
rect 304 34363 338 34397
rect 304 34295 338 34329
rect 304 34227 338 34261
rect 304 34159 338 34193
rect 304 34091 338 34125
rect 304 34023 338 34057
rect 304 33955 338 33989
rect 304 33887 338 33921
rect 304 33819 338 33853
rect 304 33751 338 33785
rect 304 33683 338 33717
rect 304 33615 338 33649
rect 304 33547 338 33581
rect 304 33479 338 33513
rect 304 33411 338 33445
rect 304 33343 338 33377
rect 304 33275 338 33309
rect 304 33207 338 33241
rect 304 33139 338 33173
rect 304 33071 338 33105
rect 304 33003 338 33037
rect 304 32935 338 32969
rect 304 32867 338 32901
rect 304 32799 338 32833
rect 304 32731 338 32765
rect 304 32663 338 32697
rect 304 32595 338 32629
rect 304 32527 338 32561
rect 304 32459 338 32493
rect 304 32391 338 32425
rect 304 32323 338 32357
rect 304 32255 338 32289
rect 304 32187 338 32221
rect 304 32119 338 32153
rect 304 32051 338 32085
rect 304 31983 338 32017
rect 304 31915 338 31949
rect 304 31847 338 31881
rect 304 31779 338 31813
rect 304 31711 338 31745
rect 304 31643 338 31677
rect 304 31575 338 31609
rect 304 31507 338 31541
rect 304 31439 338 31473
rect 304 31371 338 31405
rect 304 31303 338 31337
rect 304 31235 338 31269
rect 304 31167 338 31201
rect 304 31099 338 31133
rect 304 31031 338 31065
rect 304 30963 338 30997
rect 304 30895 338 30929
rect 304 30827 338 30861
rect 304 30759 338 30793
rect 304 30691 338 30725
rect 304 30623 338 30657
rect 304 30555 338 30589
rect 304 30487 338 30521
rect 304 30419 338 30453
rect 304 30351 338 30385
rect 304 30283 338 30317
rect 304 30215 338 30249
rect 304 30147 338 30181
rect 304 30079 338 30113
rect 304 30011 338 30045
rect 304 29943 338 29977
rect 304 29875 338 29909
rect 304 29807 338 29841
rect 304 29739 338 29773
rect 304 29671 338 29705
rect 304 29603 338 29637
rect 304 29535 338 29569
rect 304 29467 338 29501
rect 304 29399 338 29433
rect 304 29331 338 29365
rect 304 29263 338 29297
rect 304 29195 338 29229
rect 304 29127 338 29161
rect 304 29059 338 29093
rect 304 28991 338 29025
rect 304 28923 338 28957
rect 304 28855 338 28889
rect 304 28787 338 28821
rect 304 28719 338 28753
rect 304 28651 338 28685
rect 304 28583 338 28617
rect 304 28515 338 28549
rect 304 28447 338 28481
rect 304 28379 338 28413
rect 304 28311 338 28345
rect 304 28243 338 28277
rect 304 28175 338 28209
rect 304 28107 338 28141
rect 304 28039 338 28073
rect 304 27971 338 28005
rect 304 27903 338 27937
rect 304 27835 338 27869
rect 304 27767 338 27801
rect 304 27699 338 27733
rect 304 27631 338 27665
rect 304 27563 338 27597
rect 304 27495 338 27529
rect 304 27427 338 27461
rect 304 27359 338 27393
rect 304 27291 338 27325
rect 304 27223 338 27257
rect 304 27155 338 27189
rect 304 27087 338 27121
rect 304 27019 338 27053
rect 304 26951 338 26985
rect 304 26883 338 26917
rect 304 26815 338 26849
rect 304 26747 338 26781
rect 304 26679 338 26713
rect 304 26611 338 26645
rect 304 26543 338 26577
rect 304 26475 338 26509
rect 304 26407 338 26441
rect 304 26339 338 26373
rect 304 26271 338 26305
rect 304 26203 338 26237
rect 304 26135 338 26169
rect 304 26067 338 26101
rect 304 25999 338 26033
rect 304 25931 338 25965
rect 304 25863 338 25897
rect 304 25795 338 25829
rect 304 25727 338 25761
rect 304 25659 338 25693
rect 304 25591 338 25625
rect 304 25523 338 25557
rect 304 25455 338 25489
rect 304 25387 338 25421
rect 304 25319 338 25353
rect 304 25251 338 25285
rect 304 25183 338 25217
rect 304 25115 338 25149
rect 304 25047 338 25081
rect 304 24979 338 25013
rect 304 24911 338 24945
rect 304 24843 338 24877
rect 304 24775 338 24809
rect 304 24707 338 24741
rect 304 24639 338 24673
rect 304 24571 338 24605
rect 304 24503 338 24537
rect 304 24435 338 24469
rect 304 24367 338 24401
rect 304 24299 338 24333
rect 304 24231 338 24265
rect 304 24163 338 24197
rect 304 24095 338 24129
rect 304 24027 338 24061
rect 304 23959 338 23993
rect 304 23891 338 23925
rect 304 23823 338 23857
rect 304 23755 338 23789
rect 304 23687 338 23721
rect 304 23619 338 23653
rect 304 23551 338 23585
rect 304 23483 338 23517
rect 304 23415 338 23449
rect 304 23347 338 23381
rect 304 23279 338 23313
rect 304 23211 338 23245
rect 304 23143 338 23177
rect 304 23075 338 23109
rect 304 23007 338 23041
rect 304 22939 338 22973
rect 304 22871 338 22905
rect 304 22803 338 22837
rect 304 22735 338 22769
rect 304 22667 338 22701
rect 304 22599 338 22633
rect 304 22531 338 22565
rect 304 22463 338 22497
rect 304 22395 338 22429
rect 304 22327 338 22361
rect 304 22259 338 22293
rect 304 22191 338 22225
rect 304 22123 338 22157
rect 304 22055 338 22089
rect 304 21987 338 22021
rect 304 21919 338 21953
rect 304 21851 338 21885
rect 304 21783 338 21817
rect 304 21715 338 21749
rect 304 21647 338 21681
rect 304 21579 338 21613
rect 304 21511 338 21545
rect 304 21443 338 21477
rect 304 21375 338 21409
rect 304 21307 338 21341
rect 304 21239 338 21273
rect 304 21171 338 21205
rect 304 21103 338 21137
rect 304 21035 338 21069
rect 304 20967 338 21001
rect 304 20899 338 20933
rect 304 20831 338 20865
rect 304 20763 338 20797
rect 304 20695 338 20729
rect 304 20627 338 20661
rect 304 20559 338 20593
rect 304 20491 338 20525
rect 304 20423 338 20457
rect 304 20355 338 20389
rect 304 20287 338 20321
rect 304 20219 338 20253
rect 304 20151 338 20185
rect 304 20083 338 20117
rect 304 20015 338 20049
rect 304 19947 338 19981
rect 304 19879 338 19913
rect 304 19811 338 19845
rect 304 19743 338 19777
rect 304 19675 338 19709
rect 304 19607 338 19641
rect 304 19539 338 19573
rect 304 19471 338 19505
rect 304 19403 338 19437
rect 304 19335 338 19369
rect 304 19267 338 19301
rect 304 19199 338 19233
rect 304 19131 338 19165
rect 304 19063 338 19097
rect 304 18995 338 19029
rect 304 18927 338 18961
rect 304 18859 338 18893
rect 304 18791 338 18825
rect 304 18723 338 18757
rect 304 18655 338 18689
rect 304 18587 338 18621
rect 304 18519 338 18553
rect 304 18451 338 18485
rect 304 18383 338 18417
rect 304 18315 338 18349
rect 304 18247 338 18281
rect 304 18179 338 18213
rect 304 18111 338 18145
rect 304 18043 338 18077
rect 304 17975 338 18009
rect 304 17907 338 17941
rect 304 17839 338 17873
rect 304 17771 338 17805
rect 304 17703 338 17737
rect 304 17635 338 17669
rect 304 17567 338 17601
rect 304 17499 338 17533
rect 304 17431 338 17465
rect 304 17363 338 17397
rect 304 17295 338 17329
rect 304 17227 338 17261
rect 304 17159 338 17193
rect 304 17091 338 17125
rect 304 17023 338 17057
rect 304 16955 338 16989
rect 304 16887 338 16921
rect 304 16819 338 16853
rect 304 16751 338 16785
rect 304 16683 338 16717
rect 304 16615 338 16649
rect 304 16547 338 16581
rect 304 16479 338 16513
rect 304 16411 338 16445
rect 304 16343 338 16377
rect 304 16275 338 16309
rect 304 16207 338 16241
rect 304 16139 338 16173
rect 304 16071 338 16105
rect 304 16003 338 16037
rect 304 15935 338 15969
rect 304 15867 338 15901
rect 304 15799 338 15833
rect 304 15731 338 15765
rect 304 15663 338 15697
rect 304 15595 338 15629
rect 304 15527 338 15561
rect 304 15459 338 15493
rect 304 15391 338 15425
rect 304 15323 338 15357
rect 304 15255 338 15289
rect 304 15187 338 15221
rect 304 15119 338 15153
rect 304 15051 338 15085
rect 304 14983 338 15017
rect 304 14915 338 14949
rect 304 14847 338 14881
rect 304 14779 338 14813
rect 304 14711 338 14745
rect 1297 34658 1331 34692
rect 1365 34658 1399 34692
rect 1433 34658 1467 34692
rect 1501 34658 1535 34692
rect 1569 34658 1603 34692
rect 1637 34658 1671 34692
rect 1705 34658 1739 34692
rect 1773 34658 1807 34692
rect 1841 34658 1875 34692
rect 1909 34658 1943 34692
rect 1977 34658 2011 34692
rect 2045 34658 2079 34692
rect 2113 34658 2147 34692
rect 2181 34658 2215 34692
rect 2249 34658 2283 34692
rect 2317 34658 2351 34692
rect 2385 34658 2419 34692
rect 2453 34658 2487 34692
rect 2521 34658 2555 34692
rect 2589 34658 2623 34692
rect 2657 34658 2691 34692
rect 2725 34658 2759 34692
rect 2793 34658 2827 34692
rect 2861 34658 2895 34692
rect 2929 34658 2963 34692
rect 2997 34658 3031 34692
rect 3065 34658 3099 34692
rect 3133 34658 3167 34692
rect 3201 34658 3235 34692
rect 3269 34658 3303 34692
rect 3337 34658 3371 34692
rect 3405 34658 3439 34692
rect 3473 34658 3507 34692
rect 3541 34658 3575 34692
rect 3609 34658 3643 34692
rect 3677 34658 3711 34692
rect 3745 34658 3779 34692
rect 3813 34658 3847 34692
rect 3881 34658 3915 34692
rect 3949 34658 3983 34692
rect 4017 34658 4051 34692
rect 4085 34658 4119 34692
rect 4153 34658 4187 34692
rect 4221 34658 4255 34692
rect 4289 34658 4323 34692
rect 4357 34658 4391 34692
rect 4425 34658 4459 34692
rect 4493 34658 4527 34692
rect 4561 34658 4595 34692
rect 4629 34658 4663 34692
rect 4697 34658 4731 34692
rect 4765 34658 4799 34692
rect 4833 34658 4867 34692
rect 4901 34658 4935 34692
rect 4969 34658 5003 34692
rect 5037 34658 5071 34692
rect 5105 34658 5139 34692
rect 5173 34658 5207 34692
rect 5241 34658 5275 34692
rect 5309 34658 5343 34692
rect 5377 34658 5411 34692
rect 5445 34658 5479 34692
rect 5513 34658 5547 34692
rect 5581 34658 5615 34692
rect 5649 34658 5683 34692
rect 5717 34658 5751 34692
rect 5785 34658 5819 34692
rect 5853 34658 5887 34692
rect 5921 34658 5955 34692
rect 5989 34658 6023 34692
rect 6057 34658 6091 34692
rect 6125 34658 6159 34692
rect 6193 34658 6227 34692
rect 6261 34658 6295 34692
rect 6329 34658 6363 34692
rect 6397 34658 6431 34692
rect 6465 34658 6499 34692
rect 6533 34658 6567 34692
rect 6601 34658 6635 34692
rect 6669 34658 6703 34692
rect 6737 34658 6771 34692
rect 6805 34658 6839 34692
rect 6873 34658 6907 34692
rect 6941 34658 6975 34692
rect 7009 34658 7043 34692
rect 7077 34658 7111 34692
rect 7145 34658 7179 34692
rect 7213 34658 7247 34692
rect 7281 34658 7315 34692
rect 7349 34658 7383 34692
rect 7417 34658 7451 34692
rect 7485 34658 7519 34692
rect 7553 34658 7587 34692
rect 7621 34658 7655 34692
rect 7689 34658 7723 34692
rect 7757 34658 7791 34692
rect 7825 34658 7859 34692
rect 7893 34658 7927 34692
rect 7961 34658 7995 34692
rect 8029 34658 8063 34692
rect 8097 34658 8131 34692
rect 8165 34658 8199 34692
rect 8233 34658 8267 34692
rect 8301 34658 8335 34692
rect 8369 34658 8403 34692
rect 8437 34658 8471 34692
rect 8505 34658 8539 34692
rect 8573 34658 8607 34692
rect 8641 34658 8675 34692
rect 8709 34658 8743 34692
rect 8777 34658 8811 34692
rect 8845 34658 8879 34692
rect 8913 34658 8947 34692
rect 8981 34658 9015 34692
rect 9049 34658 9083 34692
rect 9117 34658 9151 34692
rect 9185 34658 9219 34692
rect 9253 34658 9287 34692
rect 9321 34658 9355 34692
rect 9389 34658 9423 34692
rect 9457 34658 9491 34692
rect 9525 34658 9559 34692
rect 9593 34658 9627 34692
rect 9661 34658 9695 34692
rect 9729 34658 9763 34692
rect 9797 34658 9831 34692
rect 9865 34658 9899 34692
rect 9933 34658 9967 34692
rect 10001 34658 10035 34692
rect 10069 34658 10103 34692
rect 10137 34658 10171 34692
rect 10205 34658 10239 34692
rect 10273 34658 10307 34692
rect 10341 34658 10375 34692
rect 10409 34658 10443 34692
rect 10477 34658 10511 34692
rect 10545 34658 10579 34692
rect 10613 34658 10647 34692
rect 10681 34658 10715 34692
rect 10749 34658 10783 34692
rect 10817 34658 10851 34692
rect 10885 34658 10919 34692
rect 10953 34658 10987 34692
rect 11021 34658 11055 34692
rect 11089 34658 11123 34692
rect 11157 34658 11191 34692
rect 11225 34658 11259 34692
rect 11293 34658 11327 34692
rect 11361 34658 11395 34692
rect 11429 34658 11463 34692
rect 11497 34658 11531 34692
rect 11565 34658 11599 34692
rect 11633 34658 11667 34692
rect 11701 34658 11735 34692
rect 11769 34658 11803 34692
rect 11837 34658 11871 34692
rect 11905 34658 11939 34692
rect 11973 34658 12007 34692
rect 12041 34658 12075 34692
rect 12109 34658 12143 34692
rect 12177 34658 12211 34692
rect 12245 34658 12279 34692
rect 12313 34658 12347 34692
rect 12381 34658 12415 34692
rect 12449 34658 12483 34692
rect 12517 34658 12551 34692
rect 12585 34658 12619 34692
rect 12653 34658 12687 34692
rect 12721 34658 12755 34692
rect 12789 34658 12823 34692
rect 12857 34658 12891 34692
rect 12925 34658 12959 34692
rect 12993 34658 13027 34692
rect 13061 34658 13095 34692
rect 13129 34658 13163 34692
rect 13197 34658 13231 34692
rect 13265 34658 13299 34692
rect 13333 34658 13367 34692
rect 13401 34658 13435 34692
rect 13469 34658 13503 34692
rect 13537 34658 13571 34692
rect 13605 34658 13639 34692
rect 13673 34658 13707 34692
rect 1153 34441 1187 34475
rect 1153 34373 1187 34407
rect 1153 34305 1187 34339
rect 1153 34237 1187 34271
rect 1153 34169 1187 34203
rect 1153 34101 1187 34135
rect 1153 34033 1187 34067
rect 1153 33965 1187 33999
rect 1153 33897 1187 33931
rect 1153 33829 1187 33863
rect 1153 33761 1187 33795
rect 1153 33693 1187 33727
rect 1153 33625 1187 33659
rect 1153 33557 1187 33591
rect 1153 33489 1187 33523
rect 1153 33421 1187 33455
rect 1153 33353 1187 33387
rect 1153 33285 1187 33319
rect 1153 33217 1187 33251
rect 1153 33149 1187 33183
rect 1153 33081 1187 33115
rect 1153 33013 1187 33047
rect 1153 32945 1187 32979
rect 1153 32877 1187 32911
rect 1153 32809 1187 32843
rect 1153 32741 1187 32775
rect 1153 32673 1187 32707
rect 1153 32605 1187 32639
rect 1153 32537 1187 32571
rect 1153 32469 1187 32503
rect 1153 32401 1187 32435
rect 1153 32333 1187 32367
rect 1153 32265 1187 32299
rect 1153 32197 1187 32231
rect 1153 32129 1187 32163
rect 1153 32061 1187 32095
rect 1153 31993 1187 32027
rect 1153 31925 1187 31959
rect 1153 31857 1187 31891
rect 1153 31789 1187 31823
rect 1153 31721 1187 31755
rect 1153 31653 1187 31687
rect 1153 31585 1187 31619
rect 1153 31517 1187 31551
rect 1153 31449 1187 31483
rect 1153 31381 1187 31415
rect 1153 31313 1187 31347
rect 1153 31245 1187 31279
rect 1153 31177 1187 31211
rect 1153 31109 1187 31143
rect 1153 31041 1187 31075
rect 1153 30973 1187 31007
rect 1153 30905 1187 30939
rect 1153 30837 1187 30871
rect 1153 30769 1187 30803
rect 1153 30701 1187 30735
rect 1153 30633 1187 30667
rect 1153 30565 1187 30599
rect 1153 30497 1187 30531
rect 1153 30429 1187 30463
rect 1153 30361 1187 30395
rect 1153 30293 1187 30327
rect 1153 30225 1187 30259
rect 1153 30157 1187 30191
rect 1153 30089 1187 30123
rect 1153 30021 1187 30055
rect 1153 29953 1187 29987
rect 1153 29885 1187 29919
rect 1153 29817 1187 29851
rect 1153 29749 1187 29783
rect 1153 29681 1187 29715
rect 1153 29613 1187 29647
rect 1153 29545 1187 29579
rect 1153 29477 1187 29511
rect 1153 29409 1187 29443
rect 1153 29341 1187 29375
rect 1153 29273 1187 29307
rect 1153 29205 1187 29239
rect 1153 29137 1187 29171
rect 1153 29069 1187 29103
rect 1153 29001 1187 29035
rect 1153 28933 1187 28967
rect 13801 34436 13835 34470
rect 13801 34368 13835 34402
rect 13801 34300 13835 34334
rect 13801 34232 13835 34266
rect 13801 34164 13835 34198
rect 13801 34096 13835 34130
rect 13801 34028 13835 34062
rect 13801 33960 13835 33994
rect 13801 33892 13835 33926
rect 13801 33824 13835 33858
rect 13801 33756 13835 33790
rect 13801 33688 13835 33722
rect 13801 33620 13835 33654
rect 13801 33552 13835 33586
rect 13801 33484 13835 33518
rect 13801 33416 13835 33450
rect 13801 33348 13835 33382
rect 13801 33280 13835 33314
rect 13801 33212 13835 33246
rect 13801 33144 13835 33178
rect 13801 33076 13835 33110
rect 13801 33008 13835 33042
rect 13801 32940 13835 32974
rect 13801 32872 13835 32906
rect 13801 32804 13835 32838
rect 13801 32736 13835 32770
rect 13801 32668 13835 32702
rect 13801 32600 13835 32634
rect 13801 32532 13835 32566
rect 13801 32464 13835 32498
rect 13801 32396 13835 32430
rect 13801 32328 13835 32362
rect 13801 32260 13835 32294
rect 13801 32192 13835 32226
rect 13801 32124 13835 32158
rect 13801 32056 13835 32090
rect 13801 31988 13835 32022
rect 13801 31920 13835 31954
rect 13801 31852 13835 31886
rect 13801 31784 13835 31818
rect 13801 31716 13835 31750
rect 13801 31648 13835 31682
rect 13801 31580 13835 31614
rect 13801 31512 13835 31546
rect 13801 31444 13835 31478
rect 13801 31376 13835 31410
rect 13801 31308 13835 31342
rect 13801 31240 13835 31274
rect 13801 31172 13835 31206
rect 13801 31104 13835 31138
rect 13801 31036 13835 31070
rect 13801 30968 13835 31002
rect 13801 30900 13835 30934
rect 13801 30832 13835 30866
rect 13801 30764 13835 30798
rect 13801 30696 13835 30730
rect 13801 30628 13835 30662
rect 13801 30560 13835 30594
rect 13801 30492 13835 30526
rect 13801 30424 13835 30458
rect 13801 30356 13835 30390
rect 13801 30288 13835 30322
rect 13801 30220 13835 30254
rect 13801 30152 13835 30186
rect 13801 30084 13835 30118
rect 13801 30016 13835 30050
rect 13801 29948 13835 29982
rect 13801 29880 13835 29914
rect 13801 29812 13835 29846
rect 13801 29744 13835 29778
rect 13801 29676 13835 29710
rect 13801 29608 13835 29642
rect 13801 29540 13835 29574
rect 13801 29472 13835 29506
rect 13801 29404 13835 29438
rect 13801 29336 13835 29370
rect 13801 29268 13835 29302
rect 13801 29200 13835 29234
rect 13801 29132 13835 29166
rect 13801 29064 13835 29098
rect 13801 28996 13835 29030
rect 13801 28928 13835 28962
rect 1153 28865 1187 28899
rect 1153 28797 1187 28831
rect 1153 28729 1187 28763
rect 1153 28661 1187 28695
rect 1153 28593 1187 28627
rect 1153 28525 1187 28559
rect 1153 28457 1187 28491
rect 1153 28389 1187 28423
rect 1153 28321 1187 28355
rect 1153 28253 1187 28287
rect 1153 28185 1187 28219
rect 1153 28117 1187 28151
rect 1153 28049 1187 28083
rect 1153 27981 1187 28015
rect 1153 27913 1187 27947
rect 1153 27845 1187 27879
rect 1153 27777 1187 27811
rect 1153 27709 1187 27743
rect 1153 27641 1187 27675
rect 1153 27573 1187 27607
rect 1153 27505 1187 27539
rect 1153 27437 1187 27471
rect 1153 27369 1187 27403
rect 1153 27301 1187 27335
rect 1153 27233 1187 27267
rect 1153 27165 1187 27199
rect 1153 27097 1187 27131
rect 1153 27029 1187 27063
rect 2485 28239 2519 28273
rect 2553 28239 2587 28273
rect 2621 28239 2655 28273
rect 2689 28239 2723 28273
rect 2757 28239 2791 28273
rect 2825 28239 2859 28273
rect 2893 28239 2927 28273
rect 2961 28239 2995 28273
rect 3029 28239 3063 28273
rect 3097 28239 3131 28273
rect 3165 28239 3199 28273
rect 3233 28239 3267 28273
rect 3301 28239 3335 28273
rect 3369 28239 3403 28273
rect 3437 28239 3471 28273
rect 3505 28239 3539 28273
rect 3573 28239 3607 28273
rect 3641 28239 3675 28273
rect 3709 28239 3743 28273
rect 3777 28239 3811 28273
rect 3845 28239 3879 28273
rect 3913 28239 3947 28273
rect 3981 28239 4015 28273
rect 4049 28239 4083 28273
rect 4117 28239 4151 28273
rect 4185 28239 4219 28273
rect 4253 28239 4287 28273
rect 4321 28239 4355 28273
rect 4389 28239 4423 28273
rect 4457 28239 4491 28273
rect 4525 28239 4559 28273
rect 4593 28239 4627 28273
rect 4661 28239 4695 28273
rect 4729 28239 4763 28273
rect 4797 28239 4831 28273
rect 4865 28239 4899 28273
rect 4933 28239 4967 28273
rect 5001 28239 5035 28273
rect 5069 28239 5103 28273
rect 5137 28239 5171 28273
rect 5205 28239 5239 28273
rect 5273 28239 5307 28273
rect 5341 28239 5375 28273
rect 5409 28239 5443 28273
rect 5477 28239 5511 28273
rect 5545 28239 5579 28273
rect 5613 28239 5647 28273
rect 5681 28239 5715 28273
rect 5749 28239 5783 28273
rect 5817 28239 5851 28273
rect 5885 28239 5919 28273
rect 5953 28239 5987 28273
rect 6021 28239 6055 28273
rect 6089 28239 6123 28273
rect 6157 28239 6191 28273
rect 6225 28239 6259 28273
rect 6293 28239 6327 28273
rect 6361 28239 6395 28273
rect 6429 28239 6463 28273
rect 6497 28239 6531 28273
rect 6565 28239 6599 28273
rect 6633 28239 6667 28273
rect 6701 28239 6735 28273
rect 6769 28239 6803 28273
rect 6837 28239 6871 28273
rect 6905 28239 6939 28273
rect 6973 28239 7007 28273
rect 7041 28239 7075 28273
rect 7109 28239 7143 28273
rect 7177 28239 7211 28273
rect 7245 28239 7279 28273
rect 7313 28239 7347 28273
rect 7381 28239 7415 28273
rect 7449 28239 7483 28273
rect 7517 28239 7551 28273
rect 7585 28239 7619 28273
rect 7653 28239 7687 28273
rect 7721 28239 7755 28273
rect 7789 28239 7823 28273
rect 7857 28239 7891 28273
rect 7925 28239 7959 28273
rect 7993 28239 8027 28273
rect 8061 28239 8095 28273
rect 8129 28239 8163 28273
rect 8197 28239 8231 28273
rect 8265 28239 8299 28273
rect 8333 28239 8367 28273
rect 8401 28239 8435 28273
rect 8469 28239 8503 28273
rect 8537 28239 8571 28273
rect 8605 28239 8639 28273
rect 8673 28239 8707 28273
rect 8741 28239 8775 28273
rect 8809 28239 8843 28273
rect 8877 28239 8911 28273
rect 8945 28239 8979 28273
rect 9013 28239 9047 28273
rect 9081 28239 9115 28273
rect 9149 28239 9183 28273
rect 9217 28239 9251 28273
rect 9285 28239 9319 28273
rect 9353 28239 9387 28273
rect 9421 28239 9455 28273
rect 9489 28239 9523 28273
rect 9557 28239 9591 28273
rect 9625 28239 9659 28273
rect 9693 28239 9727 28273
rect 9761 28239 9795 28273
rect 9829 28239 9863 28273
rect 9897 28239 9931 28273
rect 9965 28239 9999 28273
rect 10033 28239 10067 28273
rect 10101 28239 10135 28273
rect 10169 28239 10203 28273
rect 10237 28239 10271 28273
rect 10305 28239 10339 28273
rect 10373 28239 10407 28273
rect 10441 28239 10475 28273
rect 10509 28239 10543 28273
rect 10577 28239 10611 28273
rect 10645 28239 10679 28273
rect 10713 28239 10747 28273
rect 10781 28239 10815 28273
rect 10849 28239 10883 28273
rect 10917 28239 10951 28273
rect 10985 28239 11019 28273
rect 11053 28239 11087 28273
rect 11121 28239 11155 28273
rect 11189 28239 11223 28273
rect 11257 28239 11291 28273
rect 11325 28239 11359 28273
rect 11393 28239 11427 28273
rect 11461 28239 11495 28273
rect 11529 28239 11563 28273
rect 11597 28239 11631 28273
rect 11665 28239 11699 28273
rect 11733 28239 11767 28273
rect 11801 28239 11835 28273
rect 11869 28239 11903 28273
rect 11937 28239 11971 28273
rect 12005 28239 12039 28273
rect 12073 28239 12107 28273
rect 12141 28239 12175 28273
rect 12209 28239 12243 28273
rect 12277 28239 12311 28273
rect 12345 28239 12379 28273
rect 12413 28239 12447 28273
rect 12481 28239 12515 28273
rect 2485 28169 2519 28203
rect 2553 28169 2587 28203
rect 2621 28169 2655 28203
rect 2689 28169 2723 28203
rect 2757 28169 2791 28203
rect 2825 28169 2859 28203
rect 2893 28169 2927 28203
rect 2961 28169 2995 28203
rect 3029 28169 3063 28203
rect 3097 28169 3131 28203
rect 3165 28169 3199 28203
rect 3233 28169 3267 28203
rect 3301 28169 3335 28203
rect 3369 28169 3403 28203
rect 3437 28169 3471 28203
rect 3505 28169 3539 28203
rect 3573 28169 3607 28203
rect 3641 28169 3675 28203
rect 3709 28169 3743 28203
rect 3777 28169 3811 28203
rect 3845 28169 3879 28203
rect 3913 28169 3947 28203
rect 3981 28169 4015 28203
rect 4049 28169 4083 28203
rect 4117 28169 4151 28203
rect 4185 28169 4219 28203
rect 4253 28169 4287 28203
rect 4321 28169 4355 28203
rect 4389 28169 4423 28203
rect 4457 28169 4491 28203
rect 4525 28169 4559 28203
rect 4593 28169 4627 28203
rect 4661 28169 4695 28203
rect 4729 28169 4763 28203
rect 4797 28169 4831 28203
rect 4865 28169 4899 28203
rect 4933 28169 4967 28203
rect 5001 28169 5035 28203
rect 5069 28169 5103 28203
rect 5137 28169 5171 28203
rect 5205 28169 5239 28203
rect 5273 28169 5307 28203
rect 5341 28169 5375 28203
rect 5409 28169 5443 28203
rect 5477 28169 5511 28203
rect 5545 28169 5579 28203
rect 5613 28169 5647 28203
rect 5681 28169 5715 28203
rect 5749 28169 5783 28203
rect 5817 28169 5851 28203
rect 5885 28169 5919 28203
rect 5953 28169 5987 28203
rect 6021 28169 6055 28203
rect 6089 28169 6123 28203
rect 6157 28169 6191 28203
rect 6225 28169 6259 28203
rect 6293 28169 6327 28203
rect 6361 28169 6395 28203
rect 6429 28169 6463 28203
rect 6497 28169 6531 28203
rect 6565 28169 6599 28203
rect 6633 28169 6667 28203
rect 6701 28169 6735 28203
rect 6769 28169 6803 28203
rect 6837 28169 6871 28203
rect 6905 28169 6939 28203
rect 6973 28169 7007 28203
rect 7041 28169 7075 28203
rect 7109 28169 7143 28203
rect 7177 28169 7211 28203
rect 7245 28169 7279 28203
rect 7313 28169 7347 28203
rect 7381 28169 7415 28203
rect 7449 28169 7483 28203
rect 7517 28169 7551 28203
rect 7585 28169 7619 28203
rect 7653 28169 7687 28203
rect 7721 28169 7755 28203
rect 7789 28169 7823 28203
rect 7857 28169 7891 28203
rect 7925 28169 7959 28203
rect 7993 28169 8027 28203
rect 8061 28169 8095 28203
rect 8129 28169 8163 28203
rect 8197 28169 8231 28203
rect 8265 28169 8299 28203
rect 8333 28169 8367 28203
rect 8401 28169 8435 28203
rect 8469 28169 8503 28203
rect 8537 28169 8571 28203
rect 8605 28169 8639 28203
rect 8673 28169 8707 28203
rect 8741 28169 8775 28203
rect 8809 28169 8843 28203
rect 8877 28169 8911 28203
rect 8945 28169 8979 28203
rect 9013 28169 9047 28203
rect 9081 28169 9115 28203
rect 9149 28169 9183 28203
rect 9217 28169 9251 28203
rect 9285 28169 9319 28203
rect 9353 28169 9387 28203
rect 9421 28169 9455 28203
rect 9489 28169 9523 28203
rect 9557 28169 9591 28203
rect 9625 28169 9659 28203
rect 9693 28169 9727 28203
rect 9761 28169 9795 28203
rect 9829 28169 9863 28203
rect 9897 28169 9931 28203
rect 9965 28169 9999 28203
rect 10033 28169 10067 28203
rect 10101 28169 10135 28203
rect 10169 28169 10203 28203
rect 10237 28169 10271 28203
rect 10305 28169 10339 28203
rect 10373 28169 10407 28203
rect 10441 28169 10475 28203
rect 10509 28169 10543 28203
rect 10577 28169 10611 28203
rect 10645 28169 10679 28203
rect 10713 28169 10747 28203
rect 10781 28169 10815 28203
rect 10849 28169 10883 28203
rect 10917 28169 10951 28203
rect 10985 28169 11019 28203
rect 11053 28169 11087 28203
rect 11121 28169 11155 28203
rect 11189 28169 11223 28203
rect 11257 28169 11291 28203
rect 11325 28169 11359 28203
rect 11393 28169 11427 28203
rect 11461 28169 11495 28203
rect 11529 28169 11563 28203
rect 11597 28169 11631 28203
rect 11665 28169 11699 28203
rect 11733 28169 11767 28203
rect 11801 28169 11835 28203
rect 11869 28169 11903 28203
rect 11937 28169 11971 28203
rect 12005 28169 12039 28203
rect 12073 28169 12107 28203
rect 12141 28169 12175 28203
rect 12209 28169 12243 28203
rect 12277 28169 12311 28203
rect 12345 28169 12379 28203
rect 12413 28169 12447 28203
rect 12481 28169 12515 28203
rect 2376 28064 2410 28098
rect 2376 27996 2410 28030
rect 2376 27928 2410 27962
rect 2376 27860 2410 27894
rect 12590 28064 12624 28098
rect 12590 27996 12624 28030
rect 12590 27928 12624 27962
rect 12590 27860 12624 27894
rect 2485 27687 12515 27789
rect 13801 28860 13835 28894
rect 13801 28792 13835 28826
rect 13801 28724 13835 28758
rect 13801 28656 13835 28690
rect 13801 28588 13835 28622
rect 13801 28520 13835 28554
rect 13801 28452 13835 28486
rect 13801 28384 13835 28418
rect 13801 28316 13835 28350
rect 13801 28248 13835 28282
rect 13801 28180 13835 28214
rect 13801 28112 13835 28146
rect 13801 28044 13835 28078
rect 13801 27976 13835 28010
rect 13801 27908 13835 27942
rect 13801 27840 13835 27874
rect 13801 27772 13835 27806
rect 13801 27704 13835 27738
rect 13801 27636 13835 27670
rect 13801 27568 13835 27602
rect 13801 27500 13835 27534
rect 13801 27432 13835 27466
rect 13801 27364 13835 27398
rect 13801 27296 13835 27330
rect 13801 27228 13835 27262
rect 13801 27160 13835 27194
rect 13801 27092 13835 27126
rect 1153 26961 1187 26995
rect 1153 26893 1187 26927
rect 1153 26825 1187 26859
rect 1153 26757 1187 26791
rect 1153 26689 1187 26723
rect 1153 26621 1187 26655
rect 1153 26553 1187 26587
rect 13801 27024 13835 27058
rect 13801 26956 13835 26990
rect 13801 26888 13835 26922
rect 13801 26820 13835 26854
rect 13801 26752 13835 26786
rect 13801 26684 13835 26718
rect 13801 26616 13835 26650
rect 1153 26485 1187 26519
rect 1153 26417 1187 26451
rect 1153 26349 1187 26383
rect 1153 26281 1187 26315
rect 1153 26213 1187 26247
rect 1153 26145 1187 26179
rect 1153 26077 1187 26111
rect 1153 26009 1187 26043
rect 1153 25941 1187 25975
rect 1153 25873 1187 25907
rect 1153 25805 1187 25839
rect 1153 25737 1187 25771
rect 1153 25669 1187 25703
rect 1153 25601 1187 25635
rect 1153 25533 1187 25567
rect 1153 25465 1187 25499
rect 1153 25397 1187 25431
rect 1153 25329 1187 25363
rect 1153 25261 1187 25295
rect 1153 25193 1187 25227
rect 1153 25125 1187 25159
rect 1153 25057 1187 25091
rect 1153 24989 1187 25023
rect 1153 24921 1187 24955
rect 1153 24853 1187 24887
rect 2269 26201 12707 26575
rect 1758 25353 2132 26067
rect 12844 25353 13218 26067
rect 2269 24845 12707 25219
rect 13801 26548 13835 26582
rect 13801 26480 13835 26514
rect 13801 26412 13835 26446
rect 13801 26344 13835 26378
rect 13801 26276 13835 26310
rect 13801 26208 13835 26242
rect 13801 26140 13835 26174
rect 13801 26072 13835 26106
rect 13801 26004 13835 26038
rect 13801 25936 13835 25970
rect 13801 25868 13835 25902
rect 13801 25800 13835 25834
rect 13801 25732 13835 25766
rect 13801 25664 13835 25698
rect 13801 25596 13835 25630
rect 13801 25528 13835 25562
rect 13801 25460 13835 25494
rect 13801 25392 13835 25426
rect 13801 25324 13835 25358
rect 13801 25256 13835 25290
rect 13801 25188 13835 25222
rect 13801 25120 13835 25154
rect 13801 25052 13835 25086
rect 13801 24984 13835 25018
rect 13801 24916 13835 24950
rect 13801 24848 13835 24882
rect 1153 24785 1187 24819
rect 1153 24717 1187 24751
rect 1153 24649 1187 24683
rect 1153 24581 1187 24615
rect 1153 24513 1187 24547
rect 1153 24445 1187 24479
rect 1153 24377 1187 24411
rect 1153 24309 1187 24343
rect 1153 24241 1187 24275
rect 1153 24173 1187 24207
rect 1153 24105 1187 24139
rect 1153 24037 1187 24071
rect 1153 23969 1187 24003
rect 1153 23901 1187 23935
rect 1153 23833 1187 23867
rect 1153 23765 1187 23799
rect 1153 23697 1187 23731
rect 1153 23629 1187 23663
rect 1153 23561 1187 23595
rect 1153 23493 1187 23527
rect 1153 23425 1187 23459
rect 1153 23357 1187 23391
rect 1153 23289 1187 23323
rect 1153 23221 1187 23255
rect 1153 23153 1187 23187
rect 1153 23085 1187 23119
rect 1153 23017 1187 23051
rect 1153 22949 1187 22983
rect 1153 22881 1187 22915
rect 1153 22813 1187 22847
rect 1153 22745 1187 22779
rect 1153 22677 1187 22711
rect 1153 22609 1187 22643
rect 1153 22541 1187 22575
rect 1153 22473 1187 22507
rect 1153 22405 1187 22439
rect 1153 22337 1187 22371
rect 1153 22269 1187 22303
rect 1153 22201 1187 22235
rect 1153 22133 1187 22167
rect 1153 22065 1187 22099
rect 1153 21997 1187 22031
rect 1153 21929 1187 21963
rect 1153 21861 1187 21895
rect 1153 21793 1187 21827
rect 1153 21725 1187 21759
rect 1153 21657 1187 21691
rect 1153 21589 1187 21623
rect 1153 21521 1187 21555
rect 1153 21453 1187 21487
rect 1153 21385 1187 21419
rect 1153 21317 1187 21351
rect 1153 21249 1187 21283
rect 1153 21181 1187 21215
rect 1153 21113 1187 21147
rect 1153 21045 1187 21079
rect 1153 20977 1187 21011
rect 1153 20909 1187 20943
rect 1153 20841 1187 20875
rect 1153 20773 1187 20807
rect 1153 20705 1187 20739
rect 1153 20637 1187 20671
rect 1153 20569 1187 20603
rect 1153 20501 1187 20535
rect 1153 20433 1187 20467
rect 1153 20365 1187 20399
rect 1153 20297 1187 20331
rect 1153 20229 1187 20263
rect 1153 20161 1187 20195
rect 1153 20093 1187 20127
rect 1153 20025 1187 20059
rect 1153 19957 1187 19991
rect 1153 19889 1187 19923
rect 1153 19821 1187 19855
rect 1153 19753 1187 19787
rect 1153 19685 1187 19719
rect 1153 19617 1187 19651
rect 1153 19549 1187 19583
rect 1153 19481 1187 19515
rect 1153 19413 1187 19447
rect 1153 19345 1187 19379
rect 1153 19277 1187 19311
rect 1153 19209 1187 19243
rect 1153 19141 1187 19175
rect 1153 19073 1187 19107
rect 1153 19005 1187 19039
rect 1153 18937 1187 18971
rect 1153 18869 1187 18903
rect 1153 18801 1187 18835
rect 1153 18733 1187 18767
rect 1153 18665 1187 18699
rect 1153 18597 1187 18631
rect 1153 18529 1187 18563
rect 1153 18461 1187 18495
rect 1153 18393 1187 18427
rect 1153 18325 1187 18359
rect 1153 18257 1187 18291
rect 1153 18189 1187 18223
rect 1153 18121 1187 18155
rect 1153 18053 1187 18087
rect 1153 17985 1187 18019
rect 1153 17917 1187 17951
rect 1153 17849 1187 17883
rect 1153 17781 1187 17815
rect 1153 17713 1187 17747
rect 1153 17645 1187 17679
rect 1153 17577 1187 17611
rect 1153 17509 1187 17543
rect 1153 17441 1187 17475
rect 1153 17373 1187 17407
rect 1153 17305 1187 17339
rect 1153 17237 1187 17271
rect 1153 17169 1187 17203
rect 1153 17101 1187 17135
rect 1153 17033 1187 17067
rect 1153 16965 1187 16999
rect 1153 16897 1187 16931
rect 1153 16829 1187 16863
rect 1153 16761 1187 16795
rect 1153 16693 1187 16727
rect 1153 16625 1187 16659
rect 1153 16557 1187 16591
rect 1153 16489 1187 16523
rect 1153 16421 1187 16455
rect 1153 16353 1187 16387
rect 1153 16285 1187 16319
rect 1153 16217 1187 16251
rect 1153 16149 1187 16183
rect 1153 16081 1187 16115
rect 1153 16013 1187 16047
rect 1153 15945 1187 15979
rect 1153 15877 1187 15911
rect 1153 15809 1187 15843
rect 1153 15741 1187 15775
rect 1153 15673 1187 15707
rect 1153 15605 1187 15639
rect 1153 15537 1187 15571
rect 1153 15469 1187 15503
rect 1153 15401 1187 15435
rect 13801 24780 13835 24814
rect 13801 24712 13835 24746
rect 13801 24644 13835 24678
rect 13801 24576 13835 24610
rect 13801 24508 13835 24542
rect 13801 24440 13835 24474
rect 13801 24372 13835 24406
rect 13801 24304 13835 24338
rect 13801 24236 13835 24270
rect 13801 24168 13835 24202
rect 13801 24100 13835 24134
rect 13801 24032 13835 24066
rect 13801 23964 13835 23998
rect 13801 23896 13835 23930
rect 13801 23828 13835 23862
rect 13801 23760 13835 23794
rect 13801 23692 13835 23726
rect 13801 23624 13835 23658
rect 13801 23556 13835 23590
rect 13801 23488 13835 23522
rect 13801 23420 13835 23454
rect 13801 23352 13835 23386
rect 13801 23284 13835 23318
rect 13801 23216 13835 23250
rect 13801 23148 13835 23182
rect 13801 23080 13835 23114
rect 13801 23012 13835 23046
rect 13801 22944 13835 22978
rect 13801 22876 13835 22910
rect 13801 22808 13835 22842
rect 13801 22740 13835 22774
rect 13801 22672 13835 22706
rect 13801 22604 13835 22638
rect 13801 22536 13835 22570
rect 13801 22468 13835 22502
rect 13801 22400 13835 22434
rect 13801 22332 13835 22366
rect 13801 22264 13835 22298
rect 13801 22196 13835 22230
rect 13801 22128 13835 22162
rect 13801 22060 13835 22094
rect 13801 21992 13835 22026
rect 13801 21924 13835 21958
rect 13801 21856 13835 21890
rect 13801 21788 13835 21822
rect 13801 21720 13835 21754
rect 13801 21652 13835 21686
rect 13801 21584 13835 21618
rect 13801 21516 13835 21550
rect 13801 21448 13835 21482
rect 13801 21380 13835 21414
rect 13801 21312 13835 21346
rect 13801 21244 13835 21278
rect 13801 21176 13835 21210
rect 13801 21108 13835 21142
rect 13801 21040 13835 21074
rect 13801 20972 13835 21006
rect 13801 20904 13835 20938
rect 13801 20836 13835 20870
rect 13801 20768 13835 20802
rect 13801 20700 13835 20734
rect 13801 20632 13835 20666
rect 13801 20564 13835 20598
rect 13801 20496 13835 20530
rect 13801 20428 13835 20462
rect 13801 20360 13835 20394
rect 13801 20292 13835 20326
rect 13801 20224 13835 20258
rect 13801 20156 13835 20190
rect 13801 20088 13835 20122
rect 13801 20020 13835 20054
rect 13801 19952 13835 19986
rect 13801 19884 13835 19918
rect 13801 19816 13835 19850
rect 13801 19748 13835 19782
rect 13801 19680 13835 19714
rect 13801 19612 13835 19646
rect 13801 19544 13835 19578
rect 13801 19476 13835 19510
rect 13801 19408 13835 19442
rect 13801 19340 13835 19374
rect 13801 19272 13835 19306
rect 13801 19204 13835 19238
rect 13801 19136 13835 19170
rect 13801 19068 13835 19102
rect 13801 19000 13835 19034
rect 13801 18932 13835 18966
rect 13801 18864 13835 18898
rect 13801 18796 13835 18830
rect 13801 18728 13835 18762
rect 13801 18660 13835 18694
rect 13801 18592 13835 18626
rect 13801 18524 13835 18558
rect 13801 18456 13835 18490
rect 13801 18388 13835 18422
rect 13801 18320 13835 18354
rect 13801 18252 13835 18286
rect 13801 18184 13835 18218
rect 13801 18116 13835 18150
rect 13801 18048 13835 18082
rect 13801 17980 13835 18014
rect 13801 17912 13835 17946
rect 13801 17844 13835 17878
rect 13801 17776 13835 17810
rect 13801 17708 13835 17742
rect 13801 17640 13835 17674
rect 13801 17572 13835 17606
rect 13801 17504 13835 17538
rect 13801 17436 13835 17470
rect 13801 17368 13835 17402
rect 13801 17300 13835 17334
rect 13801 17232 13835 17266
rect 13801 17164 13835 17198
rect 13801 17096 13835 17130
rect 13801 17028 13835 17062
rect 13801 16960 13835 16994
rect 13801 16892 13835 16926
rect 13801 16824 13835 16858
rect 13801 16756 13835 16790
rect 13801 16688 13835 16722
rect 13801 16620 13835 16654
rect 13801 16552 13835 16586
rect 13801 16484 13835 16518
rect 13801 16416 13835 16450
rect 13801 16348 13835 16382
rect 13801 16280 13835 16314
rect 13801 16212 13835 16246
rect 13801 16144 13835 16178
rect 13801 16076 13835 16110
rect 13801 16008 13835 16042
rect 13801 15940 13835 15974
rect 13801 15872 13835 15906
rect 13801 15804 13835 15838
rect 13801 15736 13835 15770
rect 13801 15668 13835 15702
rect 13801 15600 13835 15634
rect 13801 15532 13835 15566
rect 13801 15464 13835 15498
rect 13801 15396 13835 15430
rect 1294 15257 1328 15291
rect 1362 15257 1396 15291
rect 1430 15257 1464 15291
rect 1498 15257 1532 15291
rect 1566 15257 1600 15291
rect 1634 15257 1668 15291
rect 1702 15257 1736 15291
rect 1770 15257 1804 15291
rect 1838 15257 1872 15291
rect 1906 15257 1940 15291
rect 1974 15257 2008 15291
rect 2042 15257 2076 15291
rect 2110 15257 2144 15291
rect 2178 15257 2212 15291
rect 2246 15257 2280 15291
rect 2314 15257 2348 15291
rect 2382 15257 2416 15291
rect 2450 15257 2484 15291
rect 2518 15257 2552 15291
rect 2586 15257 2620 15291
rect 2654 15257 2688 15291
rect 2722 15257 2756 15291
rect 2790 15257 2824 15291
rect 2858 15257 2892 15291
rect 2926 15257 2960 15291
rect 2994 15257 3028 15291
rect 3062 15257 3096 15291
rect 3130 15257 3164 15291
rect 3198 15257 3232 15291
rect 3266 15257 3300 15291
rect 3334 15257 3368 15291
rect 3402 15257 3436 15291
rect 3470 15257 3504 15291
rect 3538 15257 3572 15291
rect 3606 15257 3640 15291
rect 3674 15257 3708 15291
rect 3742 15257 3776 15291
rect 3810 15257 3844 15291
rect 3878 15257 3912 15291
rect 3946 15257 3980 15291
rect 4014 15257 4048 15291
rect 4082 15257 4116 15291
rect 4150 15257 4184 15291
rect 4218 15257 4252 15291
rect 4286 15257 4320 15291
rect 4354 15257 4388 15291
rect 4422 15257 4456 15291
rect 4490 15257 4524 15291
rect 4558 15257 4592 15291
rect 4626 15257 4660 15291
rect 4694 15257 4728 15291
rect 4762 15257 4796 15291
rect 4830 15257 4864 15291
rect 4898 15257 4932 15291
rect 4966 15257 5000 15291
rect 5034 15257 5068 15291
rect 5102 15257 5136 15291
rect 5170 15257 5204 15291
rect 5238 15257 5272 15291
rect 5306 15257 5340 15291
rect 5374 15257 5408 15291
rect 5442 15257 5476 15291
rect 5510 15257 5544 15291
rect 5578 15257 5612 15291
rect 5646 15257 5680 15291
rect 5714 15257 5748 15291
rect 5782 15257 5816 15291
rect 5850 15257 5884 15291
rect 5918 15257 5952 15291
rect 5986 15257 6020 15291
rect 6054 15257 6088 15291
rect 6122 15257 6156 15291
rect 6190 15257 6224 15291
rect 6258 15257 6292 15291
rect 6326 15257 6360 15291
rect 6394 15257 6428 15291
rect 6462 15257 6496 15291
rect 6530 15257 6564 15291
rect 6598 15257 6632 15291
rect 6666 15257 6700 15291
rect 6734 15257 6768 15291
rect 6802 15257 6836 15291
rect 6870 15257 6904 15291
rect 6938 15257 6972 15291
rect 7006 15257 7040 15291
rect 7074 15257 7108 15291
rect 7142 15257 7176 15291
rect 7210 15257 7244 15291
rect 7278 15257 7312 15291
rect 7346 15257 7380 15291
rect 7414 15257 7448 15291
rect 7482 15257 7516 15291
rect 7550 15257 7584 15291
rect 7618 15257 7652 15291
rect 7686 15257 7720 15291
rect 7754 15257 7788 15291
rect 7822 15257 7856 15291
rect 7890 15257 7924 15291
rect 7958 15257 7992 15291
rect 8026 15257 8060 15291
rect 8094 15257 8128 15291
rect 8162 15257 8196 15291
rect 8230 15257 8264 15291
rect 8298 15257 8332 15291
rect 8366 15257 8400 15291
rect 8434 15257 8468 15291
rect 8502 15257 8536 15291
rect 8570 15257 8604 15291
rect 8638 15257 8672 15291
rect 8706 15257 8740 15291
rect 8774 15257 8808 15291
rect 8842 15257 8876 15291
rect 8910 15257 8944 15291
rect 8978 15257 9012 15291
rect 9046 15257 9080 15291
rect 9114 15257 9148 15291
rect 9182 15257 9216 15291
rect 9250 15257 9284 15291
rect 9318 15257 9352 15291
rect 9386 15257 9420 15291
rect 9454 15257 9488 15291
rect 9522 15257 9556 15291
rect 9590 15257 9624 15291
rect 9658 15257 9692 15291
rect 9726 15257 9760 15291
rect 9794 15257 9828 15291
rect 9862 15257 9896 15291
rect 9930 15257 9964 15291
rect 9998 15257 10032 15291
rect 10066 15257 10100 15291
rect 10134 15257 10168 15291
rect 10202 15257 10236 15291
rect 10270 15257 10304 15291
rect 10338 15257 10372 15291
rect 10406 15257 10440 15291
rect 10474 15257 10508 15291
rect 10542 15257 10576 15291
rect 10610 15257 10644 15291
rect 10678 15257 10712 15291
rect 10746 15257 10780 15291
rect 10814 15257 10848 15291
rect 10882 15257 10916 15291
rect 10950 15257 10984 15291
rect 11018 15257 11052 15291
rect 11086 15257 11120 15291
rect 11154 15257 11188 15291
rect 11222 15257 11256 15291
rect 11290 15257 11324 15291
rect 11358 15257 11392 15291
rect 11426 15257 11460 15291
rect 11494 15257 11528 15291
rect 11562 15257 11596 15291
rect 11630 15257 11664 15291
rect 11698 15257 11732 15291
rect 11766 15257 11800 15291
rect 11834 15257 11868 15291
rect 11902 15257 11936 15291
rect 11970 15257 12004 15291
rect 12038 15257 12072 15291
rect 12106 15257 12140 15291
rect 12174 15257 12208 15291
rect 12242 15257 12276 15291
rect 12310 15257 12344 15291
rect 12378 15257 12412 15291
rect 12446 15257 12480 15291
rect 12514 15257 12548 15291
rect 12582 15257 12616 15291
rect 12650 15257 12684 15291
rect 12718 15257 12752 15291
rect 12786 15257 12820 15291
rect 12854 15257 12888 15291
rect 12922 15257 12956 15291
rect 12990 15257 13024 15291
rect 13058 15257 13092 15291
rect 13126 15257 13160 15291
rect 13194 15257 13228 15291
rect 13262 15257 13296 15291
rect 13330 15257 13364 15291
rect 13398 15257 13432 15291
rect 13466 15257 13500 15291
rect 13534 15257 13568 15291
rect 13602 15257 13636 15291
rect 13670 15257 13704 15291
rect 14599 36205 14633 36239
rect 14599 36137 14633 36171
rect 14599 36069 14633 36103
rect 14599 36001 14633 36035
rect 14599 35933 14633 35967
rect 14599 35865 14633 35899
rect 14599 35797 14633 35831
rect 14599 35729 14633 35763
rect 14599 35661 14633 35695
rect 14599 35593 14633 35627
rect 14599 35525 14633 35559
rect 14599 35457 14633 35491
rect 14599 35389 14633 35423
rect 14599 35321 14633 35355
rect 14599 35253 14633 35287
rect 14599 35185 14633 35219
rect 14599 35117 14633 35151
rect 14599 35049 14633 35083
rect 14599 34981 14633 35015
rect 14599 34913 14633 34947
rect 14599 34845 14633 34879
rect 14599 34777 14633 34811
rect 14599 34709 14633 34743
rect 14599 34641 14633 34675
rect 14599 34573 14633 34607
rect 14599 34505 14633 34539
rect 14599 34437 14633 34471
rect 14599 34369 14633 34403
rect 14599 34301 14633 34335
rect 14599 34233 14633 34267
rect 14599 34165 14633 34199
rect 14599 34097 14633 34131
rect 14599 34029 14633 34063
rect 14599 33961 14633 33995
rect 14599 33893 14633 33927
rect 14599 33825 14633 33859
rect 14599 33757 14633 33791
rect 14599 33689 14633 33723
rect 14599 33621 14633 33655
rect 14599 33553 14633 33587
rect 14599 33485 14633 33519
rect 14599 33417 14633 33451
rect 14599 33349 14633 33383
rect 14599 33281 14633 33315
rect 14599 33213 14633 33247
rect 14599 33145 14633 33179
rect 14599 33077 14633 33111
rect 14599 33009 14633 33043
rect 14599 32941 14633 32975
rect 14599 32873 14633 32907
rect 14599 32805 14633 32839
rect 14599 32737 14633 32771
rect 14599 32669 14633 32703
rect 14599 32601 14633 32635
rect 14599 32533 14633 32567
rect 14599 32465 14633 32499
rect 14599 32397 14633 32431
rect 14599 32329 14633 32363
rect 14599 32261 14633 32295
rect 14599 32193 14633 32227
rect 14599 32125 14633 32159
rect 14599 32057 14633 32091
rect 14599 31989 14633 32023
rect 14599 31921 14633 31955
rect 14599 31853 14633 31887
rect 14599 31785 14633 31819
rect 14599 31717 14633 31751
rect 14599 31649 14633 31683
rect 14599 31581 14633 31615
rect 14599 31513 14633 31547
rect 14599 31445 14633 31479
rect 14599 31377 14633 31411
rect 14599 31309 14633 31343
rect 14599 31241 14633 31275
rect 14599 31173 14633 31207
rect 14599 31105 14633 31139
rect 14599 31037 14633 31071
rect 14599 30969 14633 31003
rect 14599 30901 14633 30935
rect 14599 30833 14633 30867
rect 14599 30765 14633 30799
rect 14599 30697 14633 30731
rect 14599 30629 14633 30663
rect 14599 30561 14633 30595
rect 14599 30493 14633 30527
rect 14599 30425 14633 30459
rect 14599 30357 14633 30391
rect 14599 30289 14633 30323
rect 14599 30221 14633 30255
rect 14599 30153 14633 30187
rect 14599 30085 14633 30119
rect 14599 30017 14633 30051
rect 14599 29949 14633 29983
rect 14599 29881 14633 29915
rect 14599 29813 14633 29847
rect 14599 29745 14633 29779
rect 14599 29677 14633 29711
rect 14599 29609 14633 29643
rect 14599 29541 14633 29575
rect 14599 29473 14633 29507
rect 14599 29405 14633 29439
rect 14599 29337 14633 29371
rect 14599 29269 14633 29303
rect 14599 29201 14633 29235
rect 14599 29133 14633 29167
rect 14599 29065 14633 29099
rect 14599 28997 14633 29031
rect 14599 28929 14633 28963
rect 14599 28861 14633 28895
rect 14599 28793 14633 28827
rect 14599 28725 14633 28759
rect 14599 28657 14633 28691
rect 14599 28589 14633 28623
rect 14599 28521 14633 28555
rect 14599 28453 14633 28487
rect 14599 28385 14633 28419
rect 14599 28317 14633 28351
rect 14599 28249 14633 28283
rect 14599 28181 14633 28215
rect 14599 28113 14633 28147
rect 14599 28045 14633 28079
rect 14599 27977 14633 28011
rect 14599 27909 14633 27943
rect 14599 27841 14633 27875
rect 14599 27773 14633 27807
rect 14599 27705 14633 27739
rect 14599 27637 14633 27671
rect 14599 27569 14633 27603
rect 14599 27501 14633 27535
rect 14599 27433 14633 27467
rect 14599 27365 14633 27399
rect 14599 27297 14633 27331
rect 14599 27229 14633 27263
rect 14599 27161 14633 27195
rect 14599 27093 14633 27127
rect 14599 27025 14633 27059
rect 14599 26957 14633 26991
rect 14599 26889 14633 26923
rect 14599 26821 14633 26855
rect 14599 26753 14633 26787
rect 14599 26685 14633 26719
rect 14599 26617 14633 26651
rect 14599 26549 14633 26583
rect 14599 26481 14633 26515
rect 14599 26413 14633 26447
rect 14599 26345 14633 26379
rect 14599 26277 14633 26311
rect 14599 26209 14633 26243
rect 14599 26141 14633 26175
rect 14599 26073 14633 26107
rect 14599 26005 14633 26039
rect 14599 25937 14633 25971
rect 14599 25869 14633 25903
rect 14599 25801 14633 25835
rect 14599 25733 14633 25767
rect 14599 25665 14633 25699
rect 14599 25597 14633 25631
rect 14599 25529 14633 25563
rect 14599 25461 14633 25495
rect 14599 25393 14633 25427
rect 14599 25325 14633 25359
rect 14599 25257 14633 25291
rect 14599 25189 14633 25223
rect 14599 25121 14633 25155
rect 14599 25053 14633 25087
rect 14599 24985 14633 25019
rect 14599 24917 14633 24951
rect 14599 24849 14633 24883
rect 14599 24781 14633 24815
rect 14599 24713 14633 24747
rect 14599 24645 14633 24679
rect 14599 24577 14633 24611
rect 14599 24509 14633 24543
rect 14599 24441 14633 24475
rect 14599 24373 14633 24407
rect 14599 24305 14633 24339
rect 14599 24237 14633 24271
rect 14599 24169 14633 24203
rect 14599 24101 14633 24135
rect 14599 24033 14633 24067
rect 14599 23965 14633 23999
rect 14599 23897 14633 23931
rect 14599 23829 14633 23863
rect 14599 23761 14633 23795
rect 14599 23693 14633 23727
rect 14599 23625 14633 23659
rect 14599 23557 14633 23591
rect 14599 23489 14633 23523
rect 14599 23421 14633 23455
rect 14599 23353 14633 23387
rect 14599 23285 14633 23319
rect 14599 23217 14633 23251
rect 14599 23149 14633 23183
rect 14599 23081 14633 23115
rect 14599 23013 14633 23047
rect 14599 22945 14633 22979
rect 14599 22877 14633 22911
rect 14599 22809 14633 22843
rect 14599 22741 14633 22775
rect 14599 22673 14633 22707
rect 14599 22605 14633 22639
rect 14599 22537 14633 22571
rect 14599 22469 14633 22503
rect 14599 22401 14633 22435
rect 14599 22333 14633 22367
rect 14599 22265 14633 22299
rect 14599 22197 14633 22231
rect 14599 22129 14633 22163
rect 14599 22061 14633 22095
rect 14599 21993 14633 22027
rect 14599 21925 14633 21959
rect 14599 21857 14633 21891
rect 14599 21789 14633 21823
rect 14599 21721 14633 21755
rect 14599 21653 14633 21687
rect 14599 21585 14633 21619
rect 14599 21517 14633 21551
rect 14599 21449 14633 21483
rect 14599 21381 14633 21415
rect 14599 21313 14633 21347
rect 14599 21245 14633 21279
rect 14599 21177 14633 21211
rect 14599 21109 14633 21143
rect 14599 21041 14633 21075
rect 14599 20973 14633 21007
rect 14599 20905 14633 20939
rect 14599 20837 14633 20871
rect 14599 20769 14633 20803
rect 14599 20701 14633 20735
rect 14599 20633 14633 20667
rect 14599 20565 14633 20599
rect 14599 20497 14633 20531
rect 14599 20429 14633 20463
rect 14599 20361 14633 20395
rect 14599 20293 14633 20327
rect 14599 20225 14633 20259
rect 14599 20157 14633 20191
rect 14599 20089 14633 20123
rect 14599 20021 14633 20055
rect 14599 19953 14633 19987
rect 14599 19885 14633 19919
rect 14599 19817 14633 19851
rect 14599 19749 14633 19783
rect 14599 19681 14633 19715
rect 14599 19613 14633 19647
rect 14599 19545 14633 19579
rect 14599 19477 14633 19511
rect 14599 19409 14633 19443
rect 14599 19341 14633 19375
rect 14599 19273 14633 19307
rect 14599 19205 14633 19239
rect 14599 19137 14633 19171
rect 14599 19069 14633 19103
rect 14599 19001 14633 19035
rect 14599 18933 14633 18967
rect 14599 18865 14633 18899
rect 14599 18797 14633 18831
rect 14599 18729 14633 18763
rect 14599 18661 14633 18695
rect 14599 18593 14633 18627
rect 14599 18525 14633 18559
rect 14599 18457 14633 18491
rect 14599 18389 14633 18423
rect 14599 18321 14633 18355
rect 14599 18253 14633 18287
rect 14599 18185 14633 18219
rect 14599 18117 14633 18151
rect 14599 18049 14633 18083
rect 14599 17981 14633 18015
rect 14599 17913 14633 17947
rect 14599 17845 14633 17879
rect 14599 17777 14633 17811
rect 14599 17709 14633 17743
rect 14599 17641 14633 17675
rect 14599 17573 14633 17607
rect 14599 17505 14633 17539
rect 14599 17437 14633 17471
rect 14599 17369 14633 17403
rect 14599 17301 14633 17335
rect 14599 17233 14633 17267
rect 14599 17165 14633 17199
rect 14599 17097 14633 17131
rect 14599 17029 14633 17063
rect 14599 16961 14633 16995
rect 14599 16893 14633 16927
rect 14599 16825 14633 16859
rect 14599 16757 14633 16791
rect 14599 16689 14633 16723
rect 14599 16621 14633 16655
rect 14599 16553 14633 16587
rect 14599 16485 14633 16519
rect 14599 16417 14633 16451
rect 14599 16349 14633 16383
rect 14599 16281 14633 16315
rect 14599 16213 14633 16247
rect 14599 16145 14633 16179
rect 14599 16077 14633 16111
rect 14599 16009 14633 16043
rect 14599 15941 14633 15975
rect 14599 15873 14633 15907
rect 14599 15805 14633 15839
rect 14599 15737 14633 15771
rect 14599 15669 14633 15703
rect 14599 15601 14633 15635
rect 14599 15533 14633 15567
rect 14599 15465 14633 15499
rect 14599 15397 14633 15431
rect 14599 15329 14633 15363
rect 14599 15261 14633 15295
rect 14599 15193 14633 15227
rect 14599 15125 14633 15159
rect 14599 15057 14633 15091
rect 14599 14989 14633 15023
rect 14599 14921 14633 14955
rect 14599 14853 14633 14887
rect 14599 14785 14633 14819
rect 14599 14717 14633 14751
rect 304 14643 338 14677
rect 304 14575 338 14609
rect 14599 14649 14633 14683
rect 14599 14581 14633 14615
rect 468 14430 502 14464
rect 536 14430 570 14464
rect 604 14430 638 14464
rect 672 14430 706 14464
rect 740 14430 774 14464
rect 808 14430 842 14464
rect 876 14430 910 14464
rect 944 14430 978 14464
rect 1012 14430 1046 14464
rect 1080 14430 1114 14464
rect 1148 14430 1182 14464
rect 1216 14430 1250 14464
rect 1284 14430 1318 14464
rect 1352 14430 1386 14464
rect 1420 14430 1454 14464
rect 1488 14430 1522 14464
rect 1556 14430 1590 14464
rect 1624 14430 1658 14464
rect 1692 14430 1726 14464
rect 1760 14430 1794 14464
rect 1828 14430 1862 14464
rect 1896 14430 1930 14464
rect 1964 14430 1998 14464
rect 2032 14430 2066 14464
rect 2100 14430 2134 14464
rect 2168 14430 2202 14464
rect 2236 14430 2270 14464
rect 2304 14430 2338 14464
rect 2372 14430 2406 14464
rect 2440 14430 2474 14464
rect 2508 14430 2542 14464
rect 2576 14430 2610 14464
rect 2644 14430 2678 14464
rect 2712 14430 2746 14464
rect 2780 14430 2814 14464
rect 2848 14430 2882 14464
rect 2916 14430 2950 14464
rect 2984 14430 3018 14464
rect 3052 14430 3086 14464
rect 3120 14430 3154 14464
rect 3188 14430 3222 14464
rect 3256 14430 3290 14464
rect 3324 14430 3358 14464
rect 3392 14430 3426 14464
rect 3460 14430 3494 14464
rect 3528 14430 3562 14464
rect 3596 14430 3630 14464
rect 3664 14430 3698 14464
rect 3732 14430 3766 14464
rect 3800 14430 3834 14464
rect 3868 14430 3902 14464
rect 3936 14430 3970 14464
rect 4004 14430 4038 14464
rect 4072 14430 4106 14464
rect 4140 14430 4174 14464
rect 4208 14430 4242 14464
rect 4276 14430 4310 14464
rect 4344 14430 4378 14464
rect 4412 14430 4446 14464
rect 4480 14430 4514 14464
rect 4548 14430 4582 14464
rect 4616 14430 4650 14464
rect 4684 14430 4718 14464
rect 4752 14430 4786 14464
rect 4820 14430 4854 14464
rect 4888 14430 4922 14464
rect 4956 14430 4990 14464
rect 5024 14430 5058 14464
rect 5092 14430 5126 14464
rect 5160 14430 5194 14464
rect 5228 14430 5262 14464
rect 5296 14430 5330 14464
rect 5364 14430 5398 14464
rect 5432 14430 5466 14464
rect 5500 14430 5534 14464
rect 5568 14430 5602 14464
rect 5636 14430 5670 14464
rect 5704 14430 5738 14464
rect 5772 14430 5806 14464
rect 5840 14430 5874 14464
rect 5908 14430 5942 14464
rect 5976 14430 6010 14464
rect 6044 14430 6078 14464
rect 6112 14430 6146 14464
rect 6180 14430 6214 14464
rect 6248 14430 6282 14464
rect 6316 14430 6350 14464
rect 6384 14430 6418 14464
rect 6452 14430 6486 14464
rect 6520 14430 6554 14464
rect 6588 14430 6622 14464
rect 6656 14430 6690 14464
rect 6724 14430 6758 14464
rect 6792 14430 6826 14464
rect 6860 14430 6894 14464
rect 6928 14430 6962 14464
rect 6996 14430 7030 14464
rect 7064 14430 7098 14464
rect 7132 14430 7166 14464
rect 7200 14430 7234 14464
rect 7268 14430 7302 14464
rect 7336 14430 7370 14464
rect 7404 14430 7438 14464
rect 7472 14430 7506 14464
rect 7540 14430 7574 14464
rect 7608 14430 7642 14464
rect 7676 14430 7710 14464
rect 7744 14430 7778 14464
rect 7812 14430 7846 14464
rect 7880 14430 7914 14464
rect 7948 14430 7982 14464
rect 8016 14430 8050 14464
rect 8084 14430 8118 14464
rect 8152 14430 8186 14464
rect 8220 14430 8254 14464
rect 8288 14430 8322 14464
rect 8356 14430 8390 14464
rect 8424 14430 8458 14464
rect 8492 14430 8526 14464
rect 8560 14430 8594 14464
rect 8628 14430 8662 14464
rect 8696 14430 8730 14464
rect 8764 14430 8798 14464
rect 8832 14430 8866 14464
rect 8900 14430 8934 14464
rect 8968 14430 9002 14464
rect 9036 14430 9070 14464
rect 9104 14430 9138 14464
rect 9172 14430 9206 14464
rect 9240 14430 9274 14464
rect 9308 14430 9342 14464
rect 9376 14430 9410 14464
rect 9444 14430 9478 14464
rect 9512 14430 9546 14464
rect 9580 14430 9614 14464
rect 9648 14430 9682 14464
rect 9716 14430 9750 14464
rect 9784 14430 9818 14464
rect 9852 14430 9886 14464
rect 9920 14430 9954 14464
rect 9988 14430 10022 14464
rect 10056 14430 10090 14464
rect 10124 14430 10158 14464
rect 10192 14430 10226 14464
rect 10260 14430 10294 14464
rect 10328 14430 10362 14464
rect 10396 14430 10430 14464
rect 10464 14430 10498 14464
rect 10532 14430 10566 14464
rect 10600 14430 10634 14464
rect 10668 14430 10702 14464
rect 10736 14430 10770 14464
rect 10804 14430 10838 14464
rect 10872 14430 10906 14464
rect 10940 14430 10974 14464
rect 11008 14430 11042 14464
rect 11076 14430 11110 14464
rect 11144 14430 11178 14464
rect 11212 14430 11246 14464
rect 11280 14430 11314 14464
rect 11348 14430 11382 14464
rect 11416 14430 11450 14464
rect 11484 14430 11518 14464
rect 11552 14430 11586 14464
rect 11620 14430 11654 14464
rect 11688 14430 11722 14464
rect 11756 14430 11790 14464
rect 11824 14430 11858 14464
rect 11892 14430 11926 14464
rect 11960 14430 11994 14464
rect 12028 14430 12062 14464
rect 12096 14430 12130 14464
rect 12164 14430 12198 14464
rect 12232 14430 12266 14464
rect 12300 14430 12334 14464
rect 12368 14430 12402 14464
rect 12436 14430 12470 14464
rect 12504 14430 12538 14464
rect 12572 14430 12606 14464
rect 12640 14430 12674 14464
rect 12708 14430 12742 14464
rect 12776 14430 12810 14464
rect 12844 14430 12878 14464
rect 12912 14430 12946 14464
rect 12980 14430 13014 14464
rect 13048 14430 13082 14464
rect 13116 14430 13150 14464
rect 13184 14430 13218 14464
rect 13252 14430 13286 14464
rect 13320 14430 13354 14464
rect 13388 14430 13422 14464
rect 13456 14430 13490 14464
rect 13524 14430 13558 14464
rect 13592 14430 13626 14464
rect 13660 14430 13694 14464
rect 13728 14430 13762 14464
rect 13796 14430 13830 14464
rect 13864 14430 13898 14464
rect 13932 14430 13966 14464
rect 14000 14430 14034 14464
rect 14068 14430 14102 14464
rect 14136 14430 14170 14464
rect 14204 14430 14238 14464
rect 14272 14430 14306 14464
rect 14340 14430 14374 14464
rect 14408 14430 14442 14464
rect 14476 14430 14510 14464
<< mvnsubdiffcont >>
rect 758 36156 792 36190
rect 826 36156 860 36190
rect 894 36156 928 36190
rect 962 36156 996 36190
rect 1030 36156 1064 36190
rect 1098 36156 1132 36190
rect 1166 36156 1200 36190
rect 1234 36156 1268 36190
rect 1302 36156 1336 36190
rect 1370 36156 1404 36190
rect 1438 36156 1472 36190
rect 1506 36156 1540 36190
rect 1574 36156 1608 36190
rect 1642 36156 1676 36190
rect 1710 36156 1744 36190
rect 1778 36156 1812 36190
rect 1846 36156 1880 36190
rect 1914 36156 1948 36190
rect 1982 36156 2016 36190
rect 2050 36156 2084 36190
rect 2118 36156 2152 36190
rect 2186 36156 2220 36190
rect 2254 36156 2288 36190
rect 2322 36156 2356 36190
rect 2390 36156 2424 36190
rect 2458 36156 2492 36190
rect 2526 36156 2560 36190
rect 2594 36156 2628 36190
rect 2662 36156 2696 36190
rect 2730 36156 2764 36190
rect 2798 36156 2832 36190
rect 2866 36156 2900 36190
rect 2934 36156 2968 36190
rect 3002 36156 3036 36190
rect 3070 36156 3104 36190
rect 3138 36156 3172 36190
rect 3206 36156 3240 36190
rect 3274 36156 3308 36190
rect 3342 36156 3376 36190
rect 3410 36156 3444 36190
rect 3478 36156 3512 36190
rect 3546 36156 3580 36190
rect 3614 36156 3648 36190
rect 3682 36156 3716 36190
rect 3750 36156 3784 36190
rect 3818 36156 3852 36190
rect 3886 36156 3920 36190
rect 3954 36156 3988 36190
rect 4022 36156 4056 36190
rect 4090 36156 4124 36190
rect 4158 36156 4192 36190
rect 4226 36156 4260 36190
rect 4294 36156 4328 36190
rect 4362 36156 4396 36190
rect 4430 36156 4464 36190
rect 4498 36156 4532 36190
rect 4566 36156 4600 36190
rect 4634 36156 4668 36190
rect 4702 36156 4736 36190
rect 4770 36156 4804 36190
rect 4838 36156 4872 36190
rect 4906 36156 4940 36190
rect 4974 36156 5008 36190
rect 5042 36156 5076 36190
rect 5110 36156 5144 36190
rect 5178 36156 5212 36190
rect 5246 36156 5280 36190
rect 5314 36156 5348 36190
rect 5382 36156 5416 36190
rect 5450 36156 5484 36190
rect 5518 36156 5552 36190
rect 5586 36156 5620 36190
rect 5654 36156 5688 36190
rect 5722 36156 5756 36190
rect 5790 36156 5824 36190
rect 5858 36156 5892 36190
rect 5926 36156 5960 36190
rect 5994 36156 6028 36190
rect 6062 36156 6096 36190
rect 6130 36156 6164 36190
rect 6198 36156 6232 36190
rect 6266 36156 6300 36190
rect 6334 36156 6368 36190
rect 6402 36156 6436 36190
rect 6470 36156 6504 36190
rect 6538 36156 6572 36190
rect 6606 36156 6640 36190
rect 6674 36156 6708 36190
rect 6742 36156 6776 36190
rect 6810 36156 6844 36190
rect 6878 36156 6912 36190
rect 6946 36156 6980 36190
rect 7014 36156 7048 36190
rect 7082 36156 7116 36190
rect 7150 36156 7184 36190
rect 7218 36156 7252 36190
rect 7286 36156 7320 36190
rect 7354 36156 7388 36190
rect 7422 36156 7456 36190
rect 7490 36156 7524 36190
rect 7558 36156 7592 36190
rect 7626 36156 7660 36190
rect 7694 36156 7728 36190
rect 7762 36156 7796 36190
rect 7830 36156 7864 36190
rect 7898 36156 7932 36190
rect 7966 36156 8000 36190
rect 8034 36156 8068 36190
rect 8102 36156 8136 36190
rect 8170 36156 8204 36190
rect 8238 36156 8272 36190
rect 8306 36156 8340 36190
rect 8374 36156 8408 36190
rect 8442 36156 8476 36190
rect 8510 36156 8544 36190
rect 8578 36156 8612 36190
rect 8646 36156 8680 36190
rect 8714 36156 8748 36190
rect 8782 36156 8816 36190
rect 8850 36156 8884 36190
rect 8918 36156 8952 36190
rect 8986 36156 9020 36190
rect 9054 36156 9088 36190
rect 9122 36156 9156 36190
rect 9190 36156 9224 36190
rect 9258 36156 9292 36190
rect 9326 36156 9360 36190
rect 9394 36156 9428 36190
rect 9462 36156 9496 36190
rect 9530 36156 9564 36190
rect 9598 36156 9632 36190
rect 9666 36156 9700 36190
rect 9734 36156 9768 36190
rect 9802 36156 9836 36190
rect 9870 36156 9904 36190
rect 9938 36156 9972 36190
rect 10006 36156 10040 36190
rect 10074 36156 10108 36190
rect 10142 36156 10176 36190
rect 10210 36156 10244 36190
rect 10278 36156 10312 36190
rect 10346 36156 10380 36190
rect 10414 36156 10448 36190
rect 10482 36156 10516 36190
rect 10550 36156 10584 36190
rect 10618 36156 10652 36190
rect 10686 36156 10720 36190
rect 10754 36156 10788 36190
rect 10822 36156 10856 36190
rect 10890 36156 10924 36190
rect 10958 36156 10992 36190
rect 11026 36156 11060 36190
rect 11094 36156 11128 36190
rect 11162 36156 11196 36190
rect 11230 36156 11264 36190
rect 11298 36156 11332 36190
rect 11366 36156 11400 36190
rect 11434 36156 11468 36190
rect 11502 36156 11536 36190
rect 11570 36156 11604 36190
rect 11638 36156 11672 36190
rect 11706 36156 11740 36190
rect 11774 36156 11808 36190
rect 11842 36156 11876 36190
rect 11910 36156 11944 36190
rect 11978 36156 12012 36190
rect 12046 36156 12080 36190
rect 12114 36156 12148 36190
rect 12182 36156 12216 36190
rect 12250 36156 12284 36190
rect 12318 36156 12352 36190
rect 12386 36156 12420 36190
rect 12454 36156 12488 36190
rect 12522 36156 12556 36190
rect 12590 36156 12624 36190
rect 12658 36156 12692 36190
rect 12726 36156 12760 36190
rect 12794 36156 12828 36190
rect 12862 36156 12896 36190
rect 12930 36156 12964 36190
rect 12998 36156 13032 36190
rect 13066 36156 13100 36190
rect 13134 36156 13168 36190
rect 13202 36156 13236 36190
rect 13270 36156 13304 36190
rect 13338 36156 13372 36190
rect 13406 36156 13440 36190
rect 13474 36156 13508 36190
rect 13542 36156 13576 36190
rect 13610 36156 13644 36190
rect 13678 36156 13712 36190
rect 13746 36156 13780 36190
rect 13814 36156 13848 36190
rect 13882 36156 13916 36190
rect 13950 36156 13984 36190
rect 14018 36156 14052 36190
rect 14086 36156 14120 36190
rect 14154 36156 14188 36190
rect 624 36029 658 36063
rect 624 35961 658 35995
rect 624 35893 658 35927
rect 624 35825 658 35859
rect 624 35757 658 35791
rect 624 35689 658 35723
rect 624 35621 658 35655
rect 624 35553 658 35587
rect 624 35485 658 35519
rect 624 35417 658 35451
rect 624 35349 658 35383
rect 624 35281 658 35315
rect 624 35213 658 35247
rect 624 35145 658 35179
rect 624 35077 658 35111
rect 624 35009 658 35043
rect 624 34941 658 34975
rect 624 34873 658 34907
rect 624 34805 658 34839
rect 624 34737 658 34771
rect 14289 36029 14323 36063
rect 14289 35961 14323 35995
rect 14289 35893 14323 35927
rect 14289 35825 14323 35859
rect 14289 35757 14323 35791
rect 14289 35689 14323 35723
rect 14289 35621 14323 35655
rect 14289 35553 14323 35587
rect 14289 35485 14323 35519
rect 14289 35417 14323 35451
rect 14289 35349 14323 35383
rect 14289 35281 14323 35315
rect 14289 35213 14323 35247
rect 14289 35145 14323 35179
rect 14289 35077 14323 35111
rect 14289 35009 14323 35043
rect 14289 34941 14323 34975
rect 14289 34873 14323 34907
rect 14289 34805 14323 34839
rect 14289 34737 14323 34771
rect 624 34669 658 34703
rect 624 34601 658 34635
rect 624 34533 658 34567
rect 624 34465 658 34499
rect 624 34397 658 34431
rect 624 34329 658 34363
rect 624 34261 658 34295
rect 624 34193 658 34227
rect 624 34125 658 34159
rect 624 34057 658 34091
rect 624 33989 658 34023
rect 624 33921 658 33955
rect 624 33853 658 33887
rect 624 33785 658 33819
rect 624 33717 658 33751
rect 624 33649 658 33683
rect 624 33581 658 33615
rect 624 33513 658 33547
rect 624 33445 658 33479
rect 624 33377 658 33411
rect 624 33309 658 33343
rect 624 33241 658 33275
rect 624 33173 658 33207
rect 624 33105 658 33139
rect 624 33037 658 33071
rect 624 32969 658 33003
rect 624 32901 658 32935
rect 624 32833 658 32867
rect 624 32765 658 32799
rect 624 32697 658 32731
rect 624 32629 658 32663
rect 624 32561 658 32595
rect 624 32493 658 32527
rect 624 32425 658 32459
rect 624 32357 658 32391
rect 624 32289 658 32323
rect 624 32221 658 32255
rect 624 32153 658 32187
rect 624 32085 658 32119
rect 624 32017 658 32051
rect 624 31949 658 31983
rect 624 31881 658 31915
rect 624 31813 658 31847
rect 624 31745 658 31779
rect 624 31677 658 31711
rect 624 31609 658 31643
rect 624 31541 658 31575
rect 624 31473 658 31507
rect 624 31405 658 31439
rect 624 31337 658 31371
rect 624 31269 658 31303
rect 624 31201 658 31235
rect 624 31133 658 31167
rect 624 31065 658 31099
rect 624 30997 658 31031
rect 624 30929 658 30963
rect 624 30861 658 30895
rect 624 30793 658 30827
rect 624 30725 658 30759
rect 624 30657 658 30691
rect 624 30589 658 30623
rect 624 30521 658 30555
rect 624 30453 658 30487
rect 624 30385 658 30419
rect 624 30317 658 30351
rect 624 30249 658 30283
rect 624 30181 658 30215
rect 624 30113 658 30147
rect 624 30045 658 30079
rect 624 29977 658 30011
rect 624 29909 658 29943
rect 624 29841 658 29875
rect 624 29773 658 29807
rect 624 29705 658 29739
rect 624 29637 658 29671
rect 624 29569 658 29603
rect 624 29501 658 29535
rect 624 29433 658 29467
rect 624 29365 658 29399
rect 624 29297 658 29331
rect 624 29229 658 29263
rect 624 29161 658 29195
rect 624 29093 658 29127
rect 624 29025 658 29059
rect 624 28957 658 28991
rect 624 28889 658 28923
rect 624 28821 658 28855
rect 624 28753 658 28787
rect 624 28685 658 28719
rect 624 28617 658 28651
rect 624 28549 658 28583
rect 624 28481 658 28515
rect 624 28413 658 28447
rect 624 28345 658 28379
rect 624 28277 658 28311
rect 624 28209 658 28243
rect 624 28141 658 28175
rect 624 28073 658 28107
rect 624 28005 658 28039
rect 624 27937 658 27971
rect 624 27869 658 27903
rect 624 27801 658 27835
rect 624 27733 658 27767
rect 624 27665 658 27699
rect 624 27597 658 27631
rect 624 27529 658 27563
rect 624 27461 658 27495
rect 624 27393 658 27427
rect 624 27325 658 27359
rect 624 27257 658 27291
rect 624 27189 658 27223
rect 624 27121 658 27155
rect 624 27053 658 27087
rect 624 26985 658 27019
rect 624 26917 658 26951
rect 624 26849 658 26883
rect 624 26781 658 26815
rect 624 26713 658 26747
rect 624 26645 658 26679
rect 624 26577 658 26611
rect 624 26509 658 26543
rect 624 26441 658 26475
rect 624 26373 658 26407
rect 624 26305 658 26339
rect 624 26237 658 26271
rect 624 26169 658 26203
rect 624 26101 658 26135
rect 624 26033 658 26067
rect 624 25965 658 25999
rect 624 25897 658 25931
rect 624 25829 658 25863
rect 624 25761 658 25795
rect 624 25693 658 25727
rect 624 25625 658 25659
rect 624 25557 658 25591
rect 624 25489 658 25523
rect 624 25421 658 25455
rect 624 25353 658 25387
rect 624 25285 658 25319
rect 624 25217 658 25251
rect 624 25149 658 25183
rect 624 25081 658 25115
rect 624 25013 658 25047
rect 624 24945 658 24979
rect 624 24877 658 24911
rect 624 24809 658 24843
rect 624 24741 658 24775
rect 624 24673 658 24707
rect 624 24605 658 24639
rect 624 24537 658 24571
rect 624 24469 658 24503
rect 624 24401 658 24435
rect 624 24333 658 24367
rect 624 24265 658 24299
rect 624 24197 658 24231
rect 624 24129 658 24163
rect 624 24061 658 24095
rect 624 23993 658 24027
rect 624 23925 658 23959
rect 624 23857 658 23891
rect 624 23789 658 23823
rect 624 23721 658 23755
rect 624 23653 658 23687
rect 624 23585 658 23619
rect 624 23517 658 23551
rect 624 23449 658 23483
rect 624 23381 658 23415
rect 624 23313 658 23347
rect 624 23245 658 23279
rect 624 23177 658 23211
rect 624 23109 658 23143
rect 624 23041 658 23075
rect 624 22973 658 23007
rect 624 22905 658 22939
rect 624 22837 658 22871
rect 624 22769 658 22803
rect 624 22701 658 22735
rect 624 22633 658 22667
rect 624 22565 658 22599
rect 624 22497 658 22531
rect 624 22429 658 22463
rect 624 22361 658 22395
rect 624 22293 658 22327
rect 624 22225 658 22259
rect 624 22157 658 22191
rect 624 22089 658 22123
rect 624 22021 658 22055
rect 624 21953 658 21987
rect 624 21885 658 21919
rect 624 21817 658 21851
rect 624 21749 658 21783
rect 624 21681 658 21715
rect 624 21613 658 21647
rect 624 21545 658 21579
rect 624 21477 658 21511
rect 624 21409 658 21443
rect 624 21341 658 21375
rect 624 21273 658 21307
rect 624 21205 658 21239
rect 624 21137 658 21171
rect 624 21069 658 21103
rect 624 21001 658 21035
rect 624 20933 658 20967
rect 624 20865 658 20899
rect 624 20797 658 20831
rect 624 20729 658 20763
rect 624 20661 658 20695
rect 624 20593 658 20627
rect 624 20525 658 20559
rect 624 20457 658 20491
rect 624 20389 658 20423
rect 624 20321 658 20355
rect 624 20253 658 20287
rect 624 20185 658 20219
rect 624 20117 658 20151
rect 624 20049 658 20083
rect 624 19981 658 20015
rect 624 19913 658 19947
rect 624 19845 658 19879
rect 624 19777 658 19811
rect 624 19709 658 19743
rect 624 19641 658 19675
rect 624 19573 658 19607
rect 624 19505 658 19539
rect 624 19437 658 19471
rect 624 19369 658 19403
rect 624 19301 658 19335
rect 624 19233 658 19267
rect 624 19165 658 19199
rect 624 19097 658 19131
rect 624 19029 658 19063
rect 624 18961 658 18995
rect 624 18893 658 18927
rect 624 18825 658 18859
rect 624 18757 658 18791
rect 624 18689 658 18723
rect 624 18621 658 18655
rect 624 18553 658 18587
rect 624 18485 658 18519
rect 624 18417 658 18451
rect 624 18349 658 18383
rect 624 18281 658 18315
rect 624 18213 658 18247
rect 624 18145 658 18179
rect 624 18077 658 18111
rect 624 18009 658 18043
rect 624 17941 658 17975
rect 624 17873 658 17907
rect 624 17805 658 17839
rect 624 17737 658 17771
rect 624 17669 658 17703
rect 624 17601 658 17635
rect 624 17533 658 17567
rect 624 17465 658 17499
rect 624 17397 658 17431
rect 624 17329 658 17363
rect 624 17261 658 17295
rect 624 17193 658 17227
rect 624 17125 658 17159
rect 624 17057 658 17091
rect 624 16989 658 17023
rect 624 16921 658 16955
rect 624 16853 658 16887
rect 624 16785 658 16819
rect 624 16717 658 16751
rect 624 16649 658 16683
rect 624 16581 658 16615
rect 624 16513 658 16547
rect 624 16445 658 16479
rect 624 16377 658 16411
rect 624 16309 658 16343
rect 624 16241 658 16275
rect 624 16173 658 16207
rect 624 16105 658 16139
rect 624 16037 658 16071
rect 624 15969 658 16003
rect 624 15901 658 15935
rect 624 15833 658 15867
rect 624 15765 658 15799
rect 624 15697 658 15731
rect 624 15629 658 15663
rect 624 15561 658 15595
rect 624 15493 658 15527
rect 624 15425 658 15459
rect 624 15357 658 15391
rect 624 15289 658 15323
rect 624 15221 658 15255
rect 2111 28518 12889 28892
rect 1681 27517 2055 28435
rect 12945 27517 13319 28435
rect 2111 27060 12889 27434
rect 2473 25875 2507 25909
rect 2541 25875 2575 25909
rect 2609 25875 2643 25909
rect 2677 25875 2711 25909
rect 2745 25875 2779 25909
rect 2813 25875 2847 25909
rect 2881 25875 2915 25909
rect 2949 25875 2983 25909
rect 3017 25875 3051 25909
rect 3085 25875 3119 25909
rect 3153 25875 3187 25909
rect 3221 25875 3255 25909
rect 3289 25875 3323 25909
rect 3357 25875 3391 25909
rect 3425 25875 3459 25909
rect 3493 25875 3527 25909
rect 3561 25875 3595 25909
rect 3629 25875 3663 25909
rect 3697 25875 3731 25909
rect 3765 25875 3799 25909
rect 3833 25875 3867 25909
rect 3901 25875 3935 25909
rect 3969 25875 4003 25909
rect 4037 25875 4071 25909
rect 4105 25875 4139 25909
rect 4173 25875 4207 25909
rect 4241 25875 4275 25909
rect 4309 25875 4343 25909
rect 4377 25875 4411 25909
rect 4445 25875 4479 25909
rect 4513 25875 4547 25909
rect 4581 25875 4615 25909
rect 4649 25875 4683 25909
rect 4717 25875 4751 25909
rect 4785 25875 4819 25909
rect 4853 25875 4887 25909
rect 4921 25875 4955 25909
rect 4989 25875 5023 25909
rect 5057 25875 5091 25909
rect 5125 25875 5159 25909
rect 5193 25875 5227 25909
rect 5261 25875 5295 25909
rect 5329 25875 5363 25909
rect 5397 25875 5431 25909
rect 5465 25875 5499 25909
rect 5533 25875 5567 25909
rect 5601 25875 5635 25909
rect 5669 25875 5703 25909
rect 5737 25875 5771 25909
rect 5805 25875 5839 25909
rect 5873 25875 5907 25909
rect 5941 25875 5975 25909
rect 6009 25875 6043 25909
rect 6077 25875 6111 25909
rect 6145 25875 6179 25909
rect 6213 25875 6247 25909
rect 6281 25875 6315 25909
rect 6349 25875 6383 25909
rect 6417 25875 6451 25909
rect 6485 25875 6519 25909
rect 6553 25875 6587 25909
rect 6621 25875 6655 25909
rect 6689 25875 6723 25909
rect 6757 25875 6791 25909
rect 6825 25875 6859 25909
rect 6893 25875 6927 25909
rect 6961 25875 6995 25909
rect 7029 25875 7063 25909
rect 7097 25875 7131 25909
rect 7165 25875 7199 25909
rect 7233 25875 7267 25909
rect 7301 25875 7335 25909
rect 7369 25875 7403 25909
rect 7437 25875 7471 25909
rect 7505 25875 7539 25909
rect 7573 25875 7607 25909
rect 7641 25875 7675 25909
rect 7709 25875 7743 25909
rect 7777 25875 7811 25909
rect 7845 25875 7879 25909
rect 7913 25875 7947 25909
rect 7981 25875 8015 25909
rect 8049 25875 8083 25909
rect 8117 25875 8151 25909
rect 8185 25875 8219 25909
rect 8253 25875 8287 25909
rect 8321 25875 8355 25909
rect 8389 25875 8423 25909
rect 8457 25875 8491 25909
rect 8525 25875 8559 25909
rect 8593 25875 8627 25909
rect 8661 25875 8695 25909
rect 8729 25875 8763 25909
rect 8797 25875 8831 25909
rect 8865 25875 8899 25909
rect 8933 25875 8967 25909
rect 9001 25875 9035 25909
rect 9069 25875 9103 25909
rect 9137 25875 9171 25909
rect 9205 25875 9239 25909
rect 9273 25875 9307 25909
rect 9341 25875 9375 25909
rect 9409 25875 9443 25909
rect 9477 25875 9511 25909
rect 9545 25875 9579 25909
rect 9613 25875 9647 25909
rect 9681 25875 9715 25909
rect 9749 25875 9783 25909
rect 9817 25875 9851 25909
rect 9885 25875 9919 25909
rect 9953 25875 9987 25909
rect 10021 25875 10055 25909
rect 10089 25875 10123 25909
rect 10157 25875 10191 25909
rect 10225 25875 10259 25909
rect 10293 25875 10327 25909
rect 10361 25875 10395 25909
rect 10429 25875 10463 25909
rect 10497 25875 10531 25909
rect 10565 25875 10599 25909
rect 10633 25875 10667 25909
rect 10701 25875 10735 25909
rect 10769 25875 10803 25909
rect 10837 25875 10871 25909
rect 10905 25875 10939 25909
rect 10973 25875 11007 25909
rect 11041 25875 11075 25909
rect 11109 25875 11143 25909
rect 11177 25875 11211 25909
rect 11245 25875 11279 25909
rect 11313 25875 11347 25909
rect 11381 25875 11415 25909
rect 11449 25875 11483 25909
rect 11517 25875 11551 25909
rect 11585 25875 11619 25909
rect 11653 25875 11687 25909
rect 11721 25875 11755 25909
rect 11789 25875 11823 25909
rect 11857 25875 11891 25909
rect 11925 25875 11959 25909
rect 11993 25875 12027 25909
rect 12061 25875 12095 25909
rect 12129 25875 12163 25909
rect 12197 25875 12231 25909
rect 12265 25875 12299 25909
rect 12333 25875 12367 25909
rect 12401 25875 12435 25909
rect 12469 25875 12503 25909
rect 2386 25792 2420 25826
rect 2386 25724 2420 25758
rect 2386 25656 2420 25690
rect 2386 25588 2420 25622
rect 12556 25792 12590 25826
rect 12556 25724 12590 25758
rect 12556 25656 12590 25690
rect 12556 25588 12590 25622
rect 2473 25505 2507 25539
rect 2541 25505 2575 25539
rect 2609 25505 2643 25539
rect 2677 25505 2711 25539
rect 2745 25505 2779 25539
rect 2813 25505 2847 25539
rect 2881 25505 2915 25539
rect 2949 25505 2983 25539
rect 3017 25505 3051 25539
rect 3085 25505 3119 25539
rect 3153 25505 3187 25539
rect 3221 25505 3255 25539
rect 3289 25505 3323 25539
rect 3357 25505 3391 25539
rect 3425 25505 3459 25539
rect 3493 25505 3527 25539
rect 3561 25505 3595 25539
rect 3629 25505 3663 25539
rect 3697 25505 3731 25539
rect 3765 25505 3799 25539
rect 3833 25505 3867 25539
rect 3901 25505 3935 25539
rect 3969 25505 4003 25539
rect 4037 25505 4071 25539
rect 4105 25505 4139 25539
rect 4173 25505 4207 25539
rect 4241 25505 4275 25539
rect 4309 25505 4343 25539
rect 4377 25505 4411 25539
rect 4445 25505 4479 25539
rect 4513 25505 4547 25539
rect 4581 25505 4615 25539
rect 4649 25505 4683 25539
rect 4717 25505 4751 25539
rect 4785 25505 4819 25539
rect 4853 25505 4887 25539
rect 4921 25505 4955 25539
rect 4989 25505 5023 25539
rect 5057 25505 5091 25539
rect 5125 25505 5159 25539
rect 5193 25505 5227 25539
rect 5261 25505 5295 25539
rect 5329 25505 5363 25539
rect 5397 25505 5431 25539
rect 5465 25505 5499 25539
rect 5533 25505 5567 25539
rect 5601 25505 5635 25539
rect 5669 25505 5703 25539
rect 5737 25505 5771 25539
rect 5805 25505 5839 25539
rect 5873 25505 5907 25539
rect 5941 25505 5975 25539
rect 6009 25505 6043 25539
rect 6077 25505 6111 25539
rect 6145 25505 6179 25539
rect 6213 25505 6247 25539
rect 6281 25505 6315 25539
rect 6349 25505 6383 25539
rect 6417 25505 6451 25539
rect 6485 25505 6519 25539
rect 6553 25505 6587 25539
rect 6621 25505 6655 25539
rect 6689 25505 6723 25539
rect 6757 25505 6791 25539
rect 6825 25505 6859 25539
rect 6893 25505 6927 25539
rect 6961 25505 6995 25539
rect 7029 25505 7063 25539
rect 7097 25505 7131 25539
rect 7165 25505 7199 25539
rect 7233 25505 7267 25539
rect 7301 25505 7335 25539
rect 7369 25505 7403 25539
rect 7437 25505 7471 25539
rect 7505 25505 7539 25539
rect 7573 25505 7607 25539
rect 7641 25505 7675 25539
rect 7709 25505 7743 25539
rect 7777 25505 7811 25539
rect 7845 25505 7879 25539
rect 7913 25505 7947 25539
rect 7981 25505 8015 25539
rect 8049 25505 8083 25539
rect 8117 25505 8151 25539
rect 8185 25505 8219 25539
rect 8253 25505 8287 25539
rect 8321 25505 8355 25539
rect 8389 25505 8423 25539
rect 8457 25505 8491 25539
rect 8525 25505 8559 25539
rect 8593 25505 8627 25539
rect 8661 25505 8695 25539
rect 8729 25505 8763 25539
rect 8797 25505 8831 25539
rect 8865 25505 8899 25539
rect 8933 25505 8967 25539
rect 9001 25505 9035 25539
rect 9069 25505 9103 25539
rect 9137 25505 9171 25539
rect 9205 25505 9239 25539
rect 9273 25505 9307 25539
rect 9341 25505 9375 25539
rect 9409 25505 9443 25539
rect 9477 25505 9511 25539
rect 9545 25505 9579 25539
rect 9613 25505 9647 25539
rect 9681 25505 9715 25539
rect 9749 25505 9783 25539
rect 9817 25505 9851 25539
rect 9885 25505 9919 25539
rect 9953 25505 9987 25539
rect 10021 25505 10055 25539
rect 10089 25505 10123 25539
rect 10157 25505 10191 25539
rect 10225 25505 10259 25539
rect 10293 25505 10327 25539
rect 10361 25505 10395 25539
rect 10429 25505 10463 25539
rect 10497 25505 10531 25539
rect 10565 25505 10599 25539
rect 10633 25505 10667 25539
rect 10701 25505 10735 25539
rect 10769 25505 10803 25539
rect 10837 25505 10871 25539
rect 10905 25505 10939 25539
rect 10973 25505 11007 25539
rect 11041 25505 11075 25539
rect 11109 25505 11143 25539
rect 11177 25505 11211 25539
rect 11245 25505 11279 25539
rect 11313 25505 11347 25539
rect 11381 25505 11415 25539
rect 11449 25505 11483 25539
rect 11517 25505 11551 25539
rect 11585 25505 11619 25539
rect 11653 25505 11687 25539
rect 11721 25505 11755 25539
rect 11789 25505 11823 25539
rect 11857 25505 11891 25539
rect 11925 25505 11959 25539
rect 11993 25505 12027 25539
rect 12061 25505 12095 25539
rect 12129 25505 12163 25539
rect 12197 25505 12231 25539
rect 12265 25505 12299 25539
rect 12333 25505 12367 25539
rect 12401 25505 12435 25539
rect 12469 25505 12503 25539
rect 14289 34669 14323 34703
rect 14289 34601 14323 34635
rect 14289 34533 14323 34567
rect 14289 34465 14323 34499
rect 14289 34397 14323 34431
rect 14289 34329 14323 34363
rect 14289 34261 14323 34295
rect 14289 34193 14323 34227
rect 14289 34125 14323 34159
rect 14289 34057 14323 34091
rect 14289 33989 14323 34023
rect 14289 33921 14323 33955
rect 14289 33853 14323 33887
rect 14289 33785 14323 33819
rect 14289 33717 14323 33751
rect 14289 33649 14323 33683
rect 14289 33581 14323 33615
rect 14289 33513 14323 33547
rect 14289 33445 14323 33479
rect 14289 33377 14323 33411
rect 14289 33309 14323 33343
rect 14289 33241 14323 33275
rect 14289 33173 14323 33207
rect 14289 33105 14323 33139
rect 14289 33037 14323 33071
rect 14289 32969 14323 33003
rect 14289 32901 14323 32935
rect 14289 32833 14323 32867
rect 14289 32765 14323 32799
rect 14289 32697 14323 32731
rect 14289 32629 14323 32663
rect 14289 32561 14323 32595
rect 14289 32493 14323 32527
rect 14289 32425 14323 32459
rect 14289 32357 14323 32391
rect 14289 32289 14323 32323
rect 14289 32221 14323 32255
rect 14289 32153 14323 32187
rect 14289 32085 14323 32119
rect 14289 32017 14323 32051
rect 14289 31949 14323 31983
rect 14289 31881 14323 31915
rect 14289 31813 14323 31847
rect 14289 31745 14323 31779
rect 14289 31677 14323 31711
rect 14289 31609 14323 31643
rect 14289 31541 14323 31575
rect 14289 31473 14323 31507
rect 14289 31405 14323 31439
rect 14289 31337 14323 31371
rect 14289 31269 14323 31303
rect 14289 31201 14323 31235
rect 14289 31133 14323 31167
rect 14289 31065 14323 31099
rect 14289 30997 14323 31031
rect 14289 30929 14323 30963
rect 14289 30861 14323 30895
rect 14289 30793 14323 30827
rect 14289 30725 14323 30759
rect 14289 30657 14323 30691
rect 14289 30589 14323 30623
rect 14289 30521 14323 30555
rect 14289 30453 14323 30487
rect 14289 30385 14323 30419
rect 14289 30317 14323 30351
rect 14289 30249 14323 30283
rect 14289 30181 14323 30215
rect 14289 30113 14323 30147
rect 14289 30045 14323 30079
rect 14289 29977 14323 30011
rect 14289 29909 14323 29943
rect 14289 29841 14323 29875
rect 14289 29773 14323 29807
rect 14289 29705 14323 29739
rect 14289 29637 14323 29671
rect 14289 29569 14323 29603
rect 14289 29501 14323 29535
rect 14289 29433 14323 29467
rect 14289 29365 14323 29399
rect 14289 29297 14323 29331
rect 14289 29229 14323 29263
rect 14289 29161 14323 29195
rect 14289 29093 14323 29127
rect 14289 29025 14323 29059
rect 14289 28957 14323 28991
rect 14289 28889 14323 28923
rect 14289 28821 14323 28855
rect 14289 28753 14323 28787
rect 14289 28685 14323 28719
rect 14289 28617 14323 28651
rect 14289 28549 14323 28583
rect 14289 28481 14323 28515
rect 14289 28413 14323 28447
rect 14289 28345 14323 28379
rect 14289 28277 14323 28311
rect 14289 28209 14323 28243
rect 14289 28141 14323 28175
rect 14289 28073 14323 28107
rect 14289 28005 14323 28039
rect 14289 27937 14323 27971
rect 14289 27869 14323 27903
rect 14289 27801 14323 27835
rect 14289 27733 14323 27767
rect 14289 27665 14323 27699
rect 14289 27597 14323 27631
rect 14289 27529 14323 27563
rect 14289 27461 14323 27495
rect 14289 27393 14323 27427
rect 14289 27325 14323 27359
rect 14289 27257 14323 27291
rect 14289 27189 14323 27223
rect 14289 27121 14323 27155
rect 14289 27053 14323 27087
rect 14289 26985 14323 27019
rect 14289 26917 14323 26951
rect 14289 26849 14323 26883
rect 14289 26781 14323 26815
rect 14289 26713 14323 26747
rect 14289 26645 14323 26679
rect 14289 26577 14323 26611
rect 14289 26509 14323 26543
rect 14289 26441 14323 26475
rect 14289 26373 14323 26407
rect 14289 26305 14323 26339
rect 14289 26237 14323 26271
rect 14289 26169 14323 26203
rect 14289 26101 14323 26135
rect 14289 26033 14323 26067
rect 14289 25965 14323 25999
rect 14289 25897 14323 25931
rect 14289 25829 14323 25863
rect 14289 25761 14323 25795
rect 14289 25693 14323 25727
rect 14289 25625 14323 25659
rect 14289 25557 14323 25591
rect 14289 25489 14323 25523
rect 14289 25421 14323 25455
rect 14289 25353 14323 25387
rect 14289 25285 14323 25319
rect 14289 25217 14323 25251
rect 14289 25149 14323 25183
rect 14289 25081 14323 25115
rect 14289 25013 14323 25047
rect 14289 24945 14323 24979
rect 14289 24877 14323 24911
rect 14289 24809 14323 24843
rect 14289 24741 14323 24775
rect 14289 24673 14323 24707
rect 14289 24605 14323 24639
rect 14289 24537 14323 24571
rect 14289 24469 14323 24503
rect 14289 24401 14323 24435
rect 14289 24333 14323 24367
rect 14289 24265 14323 24299
rect 14289 24197 14323 24231
rect 14289 24129 14323 24163
rect 14289 24061 14323 24095
rect 14289 23993 14323 24027
rect 14289 23925 14323 23959
rect 14289 23857 14323 23891
rect 14289 23789 14323 23823
rect 14289 23721 14323 23755
rect 14289 23653 14323 23687
rect 14289 23585 14323 23619
rect 14289 23517 14323 23551
rect 14289 23449 14323 23483
rect 14289 23381 14323 23415
rect 14289 23313 14323 23347
rect 14289 23245 14323 23279
rect 14289 23177 14323 23211
rect 14289 23109 14323 23143
rect 14289 23041 14323 23075
rect 14289 22973 14323 23007
rect 14289 22905 14323 22939
rect 14289 22837 14323 22871
rect 14289 22769 14323 22803
rect 14289 22701 14323 22735
rect 14289 22633 14323 22667
rect 14289 22565 14323 22599
rect 14289 22497 14323 22531
rect 14289 22429 14323 22463
rect 14289 22361 14323 22395
rect 14289 22293 14323 22327
rect 14289 22225 14323 22259
rect 14289 22157 14323 22191
rect 14289 22089 14323 22123
rect 14289 22021 14323 22055
rect 14289 21953 14323 21987
rect 14289 21885 14323 21919
rect 14289 21817 14323 21851
rect 14289 21749 14323 21783
rect 14289 21681 14323 21715
rect 14289 21613 14323 21647
rect 14289 21545 14323 21579
rect 14289 21477 14323 21511
rect 14289 21409 14323 21443
rect 14289 21341 14323 21375
rect 14289 21273 14323 21307
rect 14289 21205 14323 21239
rect 14289 21137 14323 21171
rect 14289 21069 14323 21103
rect 14289 21001 14323 21035
rect 14289 20933 14323 20967
rect 14289 20865 14323 20899
rect 14289 20797 14323 20831
rect 14289 20729 14323 20763
rect 14289 20661 14323 20695
rect 14289 20593 14323 20627
rect 14289 20525 14323 20559
rect 14289 20457 14323 20491
rect 14289 20389 14323 20423
rect 14289 20321 14323 20355
rect 14289 20253 14323 20287
rect 14289 20185 14323 20219
rect 14289 20117 14323 20151
rect 14289 20049 14323 20083
rect 14289 19981 14323 20015
rect 14289 19913 14323 19947
rect 14289 19845 14323 19879
rect 14289 19777 14323 19811
rect 14289 19709 14323 19743
rect 14289 19641 14323 19675
rect 14289 19573 14323 19607
rect 14289 19505 14323 19539
rect 14289 19437 14323 19471
rect 14289 19369 14323 19403
rect 14289 19301 14323 19335
rect 14289 19233 14323 19267
rect 14289 19165 14323 19199
rect 14289 19097 14323 19131
rect 14289 19029 14323 19063
rect 14289 18961 14323 18995
rect 14289 18893 14323 18927
rect 14289 18825 14323 18859
rect 14289 18757 14323 18791
rect 14289 18689 14323 18723
rect 14289 18621 14323 18655
rect 14289 18553 14323 18587
rect 14289 18485 14323 18519
rect 14289 18417 14323 18451
rect 14289 18349 14323 18383
rect 14289 18281 14323 18315
rect 14289 18213 14323 18247
rect 14289 18145 14323 18179
rect 14289 18077 14323 18111
rect 14289 18009 14323 18043
rect 14289 17941 14323 17975
rect 14289 17873 14323 17907
rect 14289 17805 14323 17839
rect 14289 17737 14323 17771
rect 14289 17669 14323 17703
rect 14289 17601 14323 17635
rect 14289 17533 14323 17567
rect 14289 17465 14323 17499
rect 14289 17397 14323 17431
rect 14289 17329 14323 17363
rect 14289 17261 14323 17295
rect 14289 17193 14323 17227
rect 14289 17125 14323 17159
rect 14289 17057 14323 17091
rect 14289 16989 14323 17023
rect 14289 16921 14323 16955
rect 14289 16853 14323 16887
rect 14289 16785 14323 16819
rect 14289 16717 14323 16751
rect 14289 16649 14323 16683
rect 14289 16581 14323 16615
rect 14289 16513 14323 16547
rect 14289 16445 14323 16479
rect 14289 16377 14323 16411
rect 14289 16309 14323 16343
rect 14289 16241 14323 16275
rect 14289 16173 14323 16207
rect 14289 16105 14323 16139
rect 14289 16037 14323 16071
rect 14289 15969 14323 16003
rect 14289 15901 14323 15935
rect 14289 15833 14323 15867
rect 14289 15765 14323 15799
rect 14289 15697 14323 15731
rect 14289 15629 14323 15663
rect 14289 15561 14323 15595
rect 14289 15493 14323 15527
rect 14289 15425 14323 15459
rect 14289 15357 14323 15391
rect 14289 15289 14323 15323
rect 14289 15221 14323 15255
rect 624 15153 658 15187
rect 624 15085 658 15119
rect 624 15017 658 15051
rect 624 14949 658 14983
rect 624 14881 658 14915
rect 14289 15153 14323 15187
rect 14289 15085 14323 15119
rect 14289 15017 14323 15051
rect 14289 14949 14323 14983
rect 14289 14881 14323 14915
rect 758 14754 792 14788
rect 826 14754 860 14788
rect 894 14754 928 14788
rect 962 14754 996 14788
rect 1030 14754 1064 14788
rect 1098 14754 1132 14788
rect 1166 14754 1200 14788
rect 1234 14754 1268 14788
rect 1302 14754 1336 14788
rect 1370 14754 1404 14788
rect 1438 14754 1472 14788
rect 1506 14754 1540 14788
rect 1574 14754 1608 14788
rect 1642 14754 1676 14788
rect 1710 14754 1744 14788
rect 1778 14754 1812 14788
rect 1846 14754 1880 14788
rect 1914 14754 1948 14788
rect 1982 14754 2016 14788
rect 2050 14754 2084 14788
rect 2118 14754 2152 14788
rect 2186 14754 2220 14788
rect 2254 14754 2288 14788
rect 2322 14754 2356 14788
rect 2390 14754 2424 14788
rect 2458 14754 2492 14788
rect 2526 14754 2560 14788
rect 2594 14754 2628 14788
rect 2662 14754 2696 14788
rect 2730 14754 2764 14788
rect 2798 14754 2832 14788
rect 2866 14754 2900 14788
rect 2934 14754 2968 14788
rect 3002 14754 3036 14788
rect 3070 14754 3104 14788
rect 3138 14754 3172 14788
rect 3206 14754 3240 14788
rect 3274 14754 3308 14788
rect 3342 14754 3376 14788
rect 3410 14754 3444 14788
rect 3478 14754 3512 14788
rect 3546 14754 3580 14788
rect 3614 14754 3648 14788
rect 3682 14754 3716 14788
rect 3750 14754 3784 14788
rect 3818 14754 3852 14788
rect 3886 14754 3920 14788
rect 3954 14754 3988 14788
rect 4022 14754 4056 14788
rect 4090 14754 4124 14788
rect 4158 14754 4192 14788
rect 4226 14754 4260 14788
rect 4294 14754 4328 14788
rect 4362 14754 4396 14788
rect 4430 14754 4464 14788
rect 4498 14754 4532 14788
rect 4566 14754 4600 14788
rect 4634 14754 4668 14788
rect 4702 14754 4736 14788
rect 4770 14754 4804 14788
rect 4838 14754 4872 14788
rect 4906 14754 4940 14788
rect 4974 14754 5008 14788
rect 5042 14754 5076 14788
rect 5110 14754 5144 14788
rect 5178 14754 5212 14788
rect 5246 14754 5280 14788
rect 5314 14754 5348 14788
rect 5382 14754 5416 14788
rect 5450 14754 5484 14788
rect 5518 14754 5552 14788
rect 5586 14754 5620 14788
rect 5654 14754 5688 14788
rect 5722 14754 5756 14788
rect 5790 14754 5824 14788
rect 5858 14754 5892 14788
rect 5926 14754 5960 14788
rect 5994 14754 6028 14788
rect 6062 14754 6096 14788
rect 6130 14754 6164 14788
rect 6198 14754 6232 14788
rect 6266 14754 6300 14788
rect 6334 14754 6368 14788
rect 6402 14754 6436 14788
rect 6470 14754 6504 14788
rect 6538 14754 6572 14788
rect 6606 14754 6640 14788
rect 6674 14754 6708 14788
rect 6742 14754 6776 14788
rect 6810 14754 6844 14788
rect 6878 14754 6912 14788
rect 6946 14754 6980 14788
rect 7014 14754 7048 14788
rect 7082 14754 7116 14788
rect 7150 14754 7184 14788
rect 7218 14754 7252 14788
rect 7286 14754 7320 14788
rect 7354 14754 7388 14788
rect 7422 14754 7456 14788
rect 7490 14754 7524 14788
rect 7558 14754 7592 14788
rect 7626 14754 7660 14788
rect 7694 14754 7728 14788
rect 7762 14754 7796 14788
rect 7830 14754 7864 14788
rect 7898 14754 7932 14788
rect 7966 14754 8000 14788
rect 8034 14754 8068 14788
rect 8102 14754 8136 14788
rect 8170 14754 8204 14788
rect 8238 14754 8272 14788
rect 8306 14754 8340 14788
rect 8374 14754 8408 14788
rect 8442 14754 8476 14788
rect 8510 14754 8544 14788
rect 8578 14754 8612 14788
rect 8646 14754 8680 14788
rect 8714 14754 8748 14788
rect 8782 14754 8816 14788
rect 8850 14754 8884 14788
rect 8918 14754 8952 14788
rect 8986 14754 9020 14788
rect 9054 14754 9088 14788
rect 9122 14754 9156 14788
rect 9190 14754 9224 14788
rect 9258 14754 9292 14788
rect 9326 14754 9360 14788
rect 9394 14754 9428 14788
rect 9462 14754 9496 14788
rect 9530 14754 9564 14788
rect 9598 14754 9632 14788
rect 9666 14754 9700 14788
rect 9734 14754 9768 14788
rect 9802 14754 9836 14788
rect 9870 14754 9904 14788
rect 9938 14754 9972 14788
rect 10006 14754 10040 14788
rect 10074 14754 10108 14788
rect 10142 14754 10176 14788
rect 10210 14754 10244 14788
rect 10278 14754 10312 14788
rect 10346 14754 10380 14788
rect 10414 14754 10448 14788
rect 10482 14754 10516 14788
rect 10550 14754 10584 14788
rect 10618 14754 10652 14788
rect 10686 14754 10720 14788
rect 10754 14754 10788 14788
rect 10822 14754 10856 14788
rect 10890 14754 10924 14788
rect 10958 14754 10992 14788
rect 11026 14754 11060 14788
rect 11094 14754 11128 14788
rect 11162 14754 11196 14788
rect 11230 14754 11264 14788
rect 11298 14754 11332 14788
rect 11366 14754 11400 14788
rect 11434 14754 11468 14788
rect 11502 14754 11536 14788
rect 11570 14754 11604 14788
rect 11638 14754 11672 14788
rect 11706 14754 11740 14788
rect 11774 14754 11808 14788
rect 11842 14754 11876 14788
rect 11910 14754 11944 14788
rect 11978 14754 12012 14788
rect 12046 14754 12080 14788
rect 12114 14754 12148 14788
rect 12182 14754 12216 14788
rect 12250 14754 12284 14788
rect 12318 14754 12352 14788
rect 12386 14754 12420 14788
rect 12454 14754 12488 14788
rect 12522 14754 12556 14788
rect 12590 14754 12624 14788
rect 12658 14754 12692 14788
rect 12726 14754 12760 14788
rect 12794 14754 12828 14788
rect 12862 14754 12896 14788
rect 12930 14754 12964 14788
rect 12998 14754 13032 14788
rect 13066 14754 13100 14788
rect 13134 14754 13168 14788
rect 13202 14754 13236 14788
rect 13270 14754 13304 14788
rect 13338 14754 13372 14788
rect 13406 14754 13440 14788
rect 13474 14754 13508 14788
rect 13542 14754 13576 14788
rect 13610 14754 13644 14788
rect 13678 14754 13712 14788
rect 13746 14754 13780 14788
rect 13814 14754 13848 14788
rect 13882 14754 13916 14788
rect 13950 14754 13984 14788
rect 14018 14754 14052 14788
rect 14086 14754 14120 14788
rect 14154 14754 14188 14788
<< mvpdiode >>
rect 2488 25792 12488 25807
rect 2488 25622 2507 25792
rect 12469 25622 12488 25792
rect 2488 25607 12488 25622
<< mvndiode >>
rect 2500 28064 12500 28079
rect 2500 27894 2519 28064
rect 12481 27894 12500 28064
rect 2500 27879 12500 27894
<< mvpdiodec >>
rect 2507 25622 12469 25792
<< mvndiodec >>
rect 2519 27894 12481 28064
<< locali >>
rect 237 36547 14716 36587
rect 237 36513 312 36547
rect 346 36546 14716 36547
rect 346 36513 14606 36546
rect 237 36512 14606 36513
rect 14640 36512 14716 36546
rect 237 36511 14716 36512
rect 237 36510 548 36511
rect 582 36510 620 36511
rect 654 36510 692 36511
rect 726 36510 764 36511
rect 798 36510 836 36511
rect 870 36510 908 36511
rect 942 36510 980 36511
rect 1014 36510 1052 36511
rect 1086 36510 1124 36511
rect 1158 36510 1196 36511
rect 1230 36510 1268 36511
rect 1302 36510 1340 36511
rect 1374 36510 1412 36511
rect 1446 36510 1484 36511
rect 1518 36510 1556 36511
rect 1590 36510 1628 36511
rect 1662 36510 1700 36511
rect 1734 36510 1772 36511
rect 1806 36510 1844 36511
rect 1878 36510 1916 36511
rect 1950 36510 1988 36511
rect 2022 36510 2060 36511
rect 2094 36510 2132 36511
rect 2166 36510 2204 36511
rect 2238 36510 2276 36511
rect 2310 36510 2348 36511
rect 2382 36510 2420 36511
rect 2454 36510 2492 36511
rect 2526 36510 2564 36511
rect 2598 36510 2636 36511
rect 2670 36510 2708 36511
rect 2742 36510 2780 36511
rect 2814 36510 2852 36511
rect 2886 36510 2924 36511
rect 2958 36510 2996 36511
rect 3030 36510 3068 36511
rect 3102 36510 3140 36511
rect 3174 36510 3212 36511
rect 3246 36510 3284 36511
rect 3318 36510 3356 36511
rect 3390 36510 3428 36511
rect 3462 36510 3500 36511
rect 3534 36510 3572 36511
rect 3606 36510 3644 36511
rect 3678 36510 3716 36511
rect 3750 36510 3788 36511
rect 3822 36510 3860 36511
rect 3894 36510 3932 36511
rect 3966 36510 4004 36511
rect 4038 36510 4076 36511
rect 4110 36510 4148 36511
rect 4182 36510 4220 36511
rect 4254 36510 4292 36511
rect 4326 36510 4364 36511
rect 4398 36510 4436 36511
rect 4470 36510 4508 36511
rect 4542 36510 4580 36511
rect 4614 36510 4652 36511
rect 4686 36510 4724 36511
rect 4758 36510 4796 36511
rect 4830 36510 4868 36511
rect 4902 36510 4940 36511
rect 4974 36510 5012 36511
rect 5046 36510 5084 36511
rect 5118 36510 5156 36511
rect 5190 36510 5228 36511
rect 5262 36510 5300 36511
rect 5334 36510 5372 36511
rect 5406 36510 5444 36511
rect 5478 36510 5516 36511
rect 5550 36510 5588 36511
rect 5622 36510 5660 36511
rect 5694 36510 5732 36511
rect 5766 36510 5804 36511
rect 5838 36510 5876 36511
rect 5910 36510 5948 36511
rect 5982 36510 6020 36511
rect 6054 36510 6092 36511
rect 6126 36510 6164 36511
rect 6198 36510 6236 36511
rect 6270 36510 6308 36511
rect 6342 36510 6380 36511
rect 6414 36510 6452 36511
rect 6486 36510 6524 36511
rect 6558 36510 6596 36511
rect 6630 36510 6668 36511
rect 6702 36510 6740 36511
rect 6774 36510 6812 36511
rect 6846 36510 6884 36511
rect 6918 36510 6956 36511
rect 6990 36510 7028 36511
rect 7062 36510 7100 36511
rect 7134 36510 7172 36511
rect 7206 36510 7244 36511
rect 7278 36510 7316 36511
rect 7350 36510 7388 36511
rect 7422 36510 7460 36511
rect 7494 36510 7532 36511
rect 7566 36510 7604 36511
rect 7638 36510 7676 36511
rect 7710 36510 7748 36511
rect 7782 36510 7820 36511
rect 7854 36510 7892 36511
rect 7926 36510 7964 36511
rect 7998 36510 8036 36511
rect 8070 36510 8108 36511
rect 8142 36510 8180 36511
rect 8214 36510 8252 36511
rect 8286 36510 8324 36511
rect 8358 36510 8396 36511
rect 8430 36510 8468 36511
rect 8502 36510 8540 36511
rect 8574 36510 8612 36511
rect 8646 36510 8684 36511
rect 8718 36510 8756 36511
rect 8790 36510 8828 36511
rect 8862 36510 8900 36511
rect 8934 36510 8972 36511
rect 9006 36510 9044 36511
rect 9078 36510 9116 36511
rect 9150 36510 9188 36511
rect 9222 36510 9260 36511
rect 9294 36510 9332 36511
rect 9366 36510 9404 36511
rect 9438 36510 9476 36511
rect 9510 36510 9548 36511
rect 9582 36510 9620 36511
rect 9654 36510 9692 36511
rect 9726 36510 9764 36511
rect 9798 36510 9836 36511
rect 9870 36510 9908 36511
rect 9942 36510 9980 36511
rect 10014 36510 10052 36511
rect 10086 36510 10124 36511
rect 10158 36510 10196 36511
rect 10230 36510 10268 36511
rect 10302 36510 10340 36511
rect 10374 36510 10412 36511
rect 10446 36510 10484 36511
rect 10518 36510 10556 36511
rect 10590 36510 10628 36511
rect 10662 36510 10700 36511
rect 10734 36510 10772 36511
rect 10806 36510 10844 36511
rect 10878 36510 10916 36511
rect 10950 36510 10988 36511
rect 11022 36510 11060 36511
rect 11094 36510 11132 36511
rect 11166 36510 11204 36511
rect 11238 36510 11276 36511
rect 11310 36510 11348 36511
rect 11382 36510 11420 36511
rect 11454 36510 11492 36511
rect 11526 36510 11564 36511
rect 11598 36510 11636 36511
rect 11670 36510 11708 36511
rect 11742 36510 11780 36511
rect 11814 36510 11852 36511
rect 11886 36510 11924 36511
rect 11958 36510 11996 36511
rect 12030 36510 12068 36511
rect 12102 36510 12140 36511
rect 12174 36510 12212 36511
rect 12246 36510 12284 36511
rect 12318 36510 12356 36511
rect 12390 36510 12428 36511
rect 12462 36510 12500 36511
rect 12534 36510 12572 36511
rect 12606 36510 12644 36511
rect 12678 36510 12716 36511
rect 12750 36510 12788 36511
rect 12822 36510 12860 36511
rect 12894 36510 12932 36511
rect 12966 36510 13004 36511
rect 13038 36510 13076 36511
rect 13110 36510 13148 36511
rect 13182 36510 13220 36511
rect 13254 36510 13292 36511
rect 13326 36510 13364 36511
rect 13398 36510 13436 36511
rect 13470 36510 13508 36511
rect 13542 36510 13580 36511
rect 13614 36510 13652 36511
rect 13686 36510 13724 36511
rect 13758 36510 13796 36511
rect 13830 36510 13868 36511
rect 13902 36510 13940 36511
rect 13974 36510 14012 36511
rect 14046 36510 14084 36511
rect 14118 36510 14156 36511
rect 14190 36510 14228 36511
rect 14262 36510 14300 36511
rect 14334 36510 14372 36511
rect 14406 36510 14716 36511
rect 237 36476 447 36510
rect 481 36476 515 36510
rect 582 36477 583 36510
rect 549 36476 583 36477
rect 617 36477 620 36510
rect 685 36477 692 36510
rect 753 36477 764 36510
rect 821 36477 836 36510
rect 889 36477 908 36510
rect 957 36477 980 36510
rect 1025 36477 1052 36510
rect 1093 36477 1124 36510
rect 617 36476 651 36477
rect 685 36476 719 36477
rect 753 36476 787 36477
rect 821 36476 855 36477
rect 889 36476 923 36477
rect 957 36476 991 36477
rect 1025 36476 1059 36477
rect 1093 36476 1127 36477
rect 1161 36476 1195 36510
rect 1230 36477 1263 36510
rect 1302 36477 1331 36510
rect 1374 36477 1399 36510
rect 1446 36477 1467 36510
rect 1518 36477 1535 36510
rect 1590 36477 1603 36510
rect 1662 36477 1671 36510
rect 1734 36477 1739 36510
rect 1806 36477 1807 36510
rect 1229 36476 1263 36477
rect 1297 36476 1331 36477
rect 1365 36476 1399 36477
rect 1433 36476 1467 36477
rect 1501 36476 1535 36477
rect 1569 36476 1603 36477
rect 1637 36476 1671 36477
rect 1705 36476 1739 36477
rect 1773 36476 1807 36477
rect 1841 36477 1844 36510
rect 1909 36477 1916 36510
rect 1977 36477 1988 36510
rect 2045 36477 2060 36510
rect 2113 36477 2132 36510
rect 2181 36477 2204 36510
rect 2249 36477 2276 36510
rect 2317 36477 2348 36510
rect 1841 36476 1875 36477
rect 1909 36476 1943 36477
rect 1977 36476 2011 36477
rect 2045 36476 2079 36477
rect 2113 36476 2147 36477
rect 2181 36476 2215 36477
rect 2249 36476 2283 36477
rect 2317 36476 2351 36477
rect 2385 36476 2419 36510
rect 2454 36477 2487 36510
rect 2526 36477 2555 36510
rect 2598 36477 2623 36510
rect 2670 36477 2691 36510
rect 2742 36477 2759 36510
rect 2814 36477 2827 36510
rect 2886 36477 2895 36510
rect 2958 36477 2963 36510
rect 3030 36477 3031 36510
rect 2453 36476 2487 36477
rect 2521 36476 2555 36477
rect 2589 36476 2623 36477
rect 2657 36476 2691 36477
rect 2725 36476 2759 36477
rect 2793 36476 2827 36477
rect 2861 36476 2895 36477
rect 2929 36476 2963 36477
rect 2997 36476 3031 36477
rect 3065 36477 3068 36510
rect 3133 36477 3140 36510
rect 3201 36477 3212 36510
rect 3269 36477 3284 36510
rect 3337 36477 3356 36510
rect 3405 36477 3428 36510
rect 3473 36477 3500 36510
rect 3541 36477 3572 36510
rect 3065 36476 3099 36477
rect 3133 36476 3167 36477
rect 3201 36476 3235 36477
rect 3269 36476 3303 36477
rect 3337 36476 3371 36477
rect 3405 36476 3439 36477
rect 3473 36476 3507 36477
rect 3541 36476 3575 36477
rect 3609 36476 3643 36510
rect 3678 36477 3711 36510
rect 3750 36477 3779 36510
rect 3822 36477 3847 36510
rect 3894 36477 3915 36510
rect 3966 36477 3983 36510
rect 4038 36477 4051 36510
rect 4110 36477 4119 36510
rect 4182 36477 4187 36510
rect 4254 36477 4255 36510
rect 3677 36476 3711 36477
rect 3745 36476 3779 36477
rect 3813 36476 3847 36477
rect 3881 36476 3915 36477
rect 3949 36476 3983 36477
rect 4017 36476 4051 36477
rect 4085 36476 4119 36477
rect 4153 36476 4187 36477
rect 4221 36476 4255 36477
rect 4289 36477 4292 36510
rect 4357 36477 4364 36510
rect 4425 36477 4436 36510
rect 4493 36477 4508 36510
rect 4561 36477 4580 36510
rect 4629 36477 4652 36510
rect 4697 36477 4724 36510
rect 4765 36477 4796 36510
rect 4289 36476 4323 36477
rect 4357 36476 4391 36477
rect 4425 36476 4459 36477
rect 4493 36476 4527 36477
rect 4561 36476 4595 36477
rect 4629 36476 4663 36477
rect 4697 36476 4731 36477
rect 4765 36476 4799 36477
rect 4833 36476 4867 36510
rect 4902 36477 4935 36510
rect 4974 36477 5003 36510
rect 5046 36477 5071 36510
rect 5118 36477 5139 36510
rect 5190 36477 5207 36510
rect 5262 36477 5275 36510
rect 5334 36477 5343 36510
rect 5406 36477 5411 36510
rect 5478 36477 5479 36510
rect 4901 36476 4935 36477
rect 4969 36476 5003 36477
rect 5037 36476 5071 36477
rect 5105 36476 5139 36477
rect 5173 36476 5207 36477
rect 5241 36476 5275 36477
rect 5309 36476 5343 36477
rect 5377 36476 5411 36477
rect 5445 36476 5479 36477
rect 5513 36477 5516 36510
rect 5581 36477 5588 36510
rect 5649 36477 5660 36510
rect 5717 36477 5732 36510
rect 5785 36477 5804 36510
rect 5853 36477 5876 36510
rect 5921 36477 5948 36510
rect 5989 36477 6020 36510
rect 5513 36476 5547 36477
rect 5581 36476 5615 36477
rect 5649 36476 5683 36477
rect 5717 36476 5751 36477
rect 5785 36476 5819 36477
rect 5853 36476 5887 36477
rect 5921 36476 5955 36477
rect 5989 36476 6023 36477
rect 6057 36476 6091 36510
rect 6126 36477 6159 36510
rect 6198 36477 6227 36510
rect 6270 36477 6295 36510
rect 6342 36477 6363 36510
rect 6414 36477 6431 36510
rect 6486 36477 6499 36510
rect 6558 36477 6567 36510
rect 6630 36477 6635 36510
rect 6702 36477 6703 36510
rect 6125 36476 6159 36477
rect 6193 36476 6227 36477
rect 6261 36476 6295 36477
rect 6329 36476 6363 36477
rect 6397 36476 6431 36477
rect 6465 36476 6499 36477
rect 6533 36476 6567 36477
rect 6601 36476 6635 36477
rect 6669 36476 6703 36477
rect 6737 36477 6740 36510
rect 6805 36477 6812 36510
rect 6873 36477 6884 36510
rect 6941 36477 6956 36510
rect 7009 36477 7028 36510
rect 7077 36477 7100 36510
rect 7145 36477 7172 36510
rect 7213 36477 7244 36510
rect 6737 36476 6771 36477
rect 6805 36476 6839 36477
rect 6873 36476 6907 36477
rect 6941 36476 6975 36477
rect 7009 36476 7043 36477
rect 7077 36476 7111 36477
rect 7145 36476 7179 36477
rect 7213 36476 7247 36477
rect 7281 36476 7315 36510
rect 7350 36477 7383 36510
rect 7422 36477 7451 36510
rect 7494 36477 7519 36510
rect 7566 36477 7587 36510
rect 7638 36477 7655 36510
rect 7710 36477 7723 36510
rect 7782 36477 7791 36510
rect 7854 36477 7859 36510
rect 7926 36477 7927 36510
rect 7349 36476 7383 36477
rect 7417 36476 7451 36477
rect 7485 36476 7519 36477
rect 7553 36476 7587 36477
rect 7621 36476 7655 36477
rect 7689 36476 7723 36477
rect 7757 36476 7791 36477
rect 7825 36476 7859 36477
rect 7893 36476 7927 36477
rect 7961 36477 7964 36510
rect 8029 36477 8036 36510
rect 8097 36477 8108 36510
rect 8165 36477 8180 36510
rect 8233 36477 8252 36510
rect 8301 36477 8324 36510
rect 8369 36477 8396 36510
rect 8437 36477 8468 36510
rect 7961 36476 7995 36477
rect 8029 36476 8063 36477
rect 8097 36476 8131 36477
rect 8165 36476 8199 36477
rect 8233 36476 8267 36477
rect 8301 36476 8335 36477
rect 8369 36476 8403 36477
rect 8437 36476 8471 36477
rect 8505 36476 8539 36510
rect 8574 36477 8607 36510
rect 8646 36477 8675 36510
rect 8718 36477 8743 36510
rect 8790 36477 8811 36510
rect 8862 36477 8879 36510
rect 8934 36477 8947 36510
rect 9006 36477 9015 36510
rect 9078 36477 9083 36510
rect 9150 36477 9151 36510
rect 8573 36476 8607 36477
rect 8641 36476 8675 36477
rect 8709 36476 8743 36477
rect 8777 36476 8811 36477
rect 8845 36476 8879 36477
rect 8913 36476 8947 36477
rect 8981 36476 9015 36477
rect 9049 36476 9083 36477
rect 9117 36476 9151 36477
rect 9185 36477 9188 36510
rect 9253 36477 9260 36510
rect 9321 36477 9332 36510
rect 9389 36477 9404 36510
rect 9457 36477 9476 36510
rect 9525 36477 9548 36510
rect 9593 36477 9620 36510
rect 9661 36477 9692 36510
rect 9185 36476 9219 36477
rect 9253 36476 9287 36477
rect 9321 36476 9355 36477
rect 9389 36476 9423 36477
rect 9457 36476 9491 36477
rect 9525 36476 9559 36477
rect 9593 36476 9627 36477
rect 9661 36476 9695 36477
rect 9729 36476 9763 36510
rect 9798 36477 9831 36510
rect 9870 36477 9899 36510
rect 9942 36477 9967 36510
rect 10014 36477 10035 36510
rect 10086 36477 10103 36510
rect 10158 36477 10171 36510
rect 10230 36477 10239 36510
rect 10302 36477 10307 36510
rect 10374 36477 10375 36510
rect 9797 36476 9831 36477
rect 9865 36476 9899 36477
rect 9933 36476 9967 36477
rect 10001 36476 10035 36477
rect 10069 36476 10103 36477
rect 10137 36476 10171 36477
rect 10205 36476 10239 36477
rect 10273 36476 10307 36477
rect 10341 36476 10375 36477
rect 10409 36477 10412 36510
rect 10477 36477 10484 36510
rect 10545 36477 10556 36510
rect 10613 36477 10628 36510
rect 10681 36477 10700 36510
rect 10749 36477 10772 36510
rect 10817 36477 10844 36510
rect 10885 36477 10916 36510
rect 10409 36476 10443 36477
rect 10477 36476 10511 36477
rect 10545 36476 10579 36477
rect 10613 36476 10647 36477
rect 10681 36476 10715 36477
rect 10749 36476 10783 36477
rect 10817 36476 10851 36477
rect 10885 36476 10919 36477
rect 10953 36476 10987 36510
rect 11022 36477 11055 36510
rect 11094 36477 11123 36510
rect 11166 36477 11191 36510
rect 11238 36477 11259 36510
rect 11310 36477 11327 36510
rect 11382 36477 11395 36510
rect 11454 36477 11463 36510
rect 11526 36477 11531 36510
rect 11598 36477 11599 36510
rect 11021 36476 11055 36477
rect 11089 36476 11123 36477
rect 11157 36476 11191 36477
rect 11225 36476 11259 36477
rect 11293 36476 11327 36477
rect 11361 36476 11395 36477
rect 11429 36476 11463 36477
rect 11497 36476 11531 36477
rect 11565 36476 11599 36477
rect 11633 36477 11636 36510
rect 11701 36477 11708 36510
rect 11769 36477 11780 36510
rect 11837 36477 11852 36510
rect 11905 36477 11924 36510
rect 11973 36477 11996 36510
rect 12041 36477 12068 36510
rect 12109 36477 12140 36510
rect 11633 36476 11667 36477
rect 11701 36476 11735 36477
rect 11769 36476 11803 36477
rect 11837 36476 11871 36477
rect 11905 36476 11939 36477
rect 11973 36476 12007 36477
rect 12041 36476 12075 36477
rect 12109 36476 12143 36477
rect 12177 36476 12211 36510
rect 12246 36477 12279 36510
rect 12318 36477 12347 36510
rect 12390 36477 12415 36510
rect 12462 36477 12483 36510
rect 12534 36477 12551 36510
rect 12606 36477 12619 36510
rect 12678 36477 12687 36510
rect 12750 36477 12755 36510
rect 12822 36477 12823 36510
rect 12245 36476 12279 36477
rect 12313 36476 12347 36477
rect 12381 36476 12415 36477
rect 12449 36476 12483 36477
rect 12517 36476 12551 36477
rect 12585 36476 12619 36477
rect 12653 36476 12687 36477
rect 12721 36476 12755 36477
rect 12789 36476 12823 36477
rect 12857 36477 12860 36510
rect 12925 36477 12932 36510
rect 12993 36477 13004 36510
rect 13061 36477 13076 36510
rect 13129 36477 13148 36510
rect 13197 36477 13220 36510
rect 13265 36477 13292 36510
rect 13333 36477 13364 36510
rect 12857 36476 12891 36477
rect 12925 36476 12959 36477
rect 12993 36476 13027 36477
rect 13061 36476 13095 36477
rect 13129 36476 13163 36477
rect 13197 36476 13231 36477
rect 13265 36476 13299 36477
rect 13333 36476 13367 36477
rect 13401 36476 13435 36510
rect 13470 36477 13503 36510
rect 13542 36477 13571 36510
rect 13614 36477 13639 36510
rect 13686 36477 13707 36510
rect 13758 36477 13775 36510
rect 13830 36477 13843 36510
rect 13902 36477 13911 36510
rect 13974 36477 13979 36510
rect 14046 36477 14047 36510
rect 13469 36476 13503 36477
rect 13537 36476 13571 36477
rect 13605 36476 13639 36477
rect 13673 36476 13707 36477
rect 13741 36476 13775 36477
rect 13809 36476 13843 36477
rect 13877 36476 13911 36477
rect 13945 36476 13979 36477
rect 14013 36476 14047 36477
rect 14081 36477 14084 36510
rect 14149 36477 14156 36510
rect 14217 36477 14228 36510
rect 14285 36477 14300 36510
rect 14353 36477 14372 36510
rect 14081 36476 14115 36477
rect 14149 36476 14183 36477
rect 14217 36476 14251 36477
rect 14285 36476 14319 36477
rect 14353 36476 14387 36477
rect 14421 36476 14455 36510
rect 14489 36476 14716 36510
rect 237 36475 14716 36476
rect 237 36441 312 36475
rect 346 36474 14716 36475
rect 346 36441 14606 36474
rect 237 36440 14606 36441
rect 14640 36440 14716 36474
rect 237 36402 14716 36440
rect 237 36369 422 36402
rect 237 36335 304 36369
rect 338 36335 422 36369
rect 237 36301 422 36335
rect 237 36267 304 36301
rect 338 36294 422 36301
rect 237 36260 312 36267
rect 346 36260 422 36294
rect 237 36233 422 36260
rect 237 36199 304 36233
rect 338 36222 422 36233
rect 237 36188 312 36199
rect 346 36188 422 36222
rect 14531 36375 14716 36402
rect 14531 36341 14599 36375
rect 14633 36341 14716 36375
rect 14531 36307 14716 36341
rect 14531 36273 14599 36307
rect 14633 36291 14716 36307
rect 14531 36257 14606 36273
rect 14640 36257 14716 36291
rect 14531 36239 14716 36257
rect 237 36165 422 36188
rect 237 36131 304 36165
rect 338 36150 422 36165
rect 237 36116 312 36131
rect 346 36116 422 36150
rect 237 36097 422 36116
rect 237 36063 304 36097
rect 338 36078 422 36097
rect 237 36044 312 36063
rect 346 36044 422 36078
rect 237 36029 422 36044
rect 237 35995 304 36029
rect 338 36006 422 36029
rect 237 35972 312 35995
rect 346 35972 422 36006
rect 237 35961 422 35972
rect 237 35927 304 35961
rect 338 35934 422 35961
rect 237 35900 312 35927
rect 346 35900 422 35934
rect 237 35893 422 35900
rect 237 35859 304 35893
rect 338 35862 422 35893
rect 237 35828 312 35859
rect 346 35828 422 35862
rect 237 35825 422 35828
rect 237 35791 304 35825
rect 338 35791 422 35825
rect 237 35790 422 35791
rect 237 35757 312 35790
rect 237 35723 304 35757
rect 346 35756 422 35790
rect 338 35723 422 35756
rect 237 35718 422 35723
rect 237 35689 312 35718
rect 237 35655 304 35689
rect 346 35684 422 35718
rect 338 35655 422 35684
rect 237 35646 422 35655
rect 237 35621 312 35646
rect 237 35587 304 35621
rect 346 35612 422 35646
rect 338 35587 422 35612
rect 237 35574 422 35587
rect 237 35553 312 35574
rect 237 35519 304 35553
rect 346 35540 422 35574
rect 338 35519 422 35540
rect 237 35502 422 35519
rect 237 35485 312 35502
rect 237 35451 304 35485
rect 346 35468 422 35502
rect 338 35451 422 35468
rect 237 35430 422 35451
rect 237 35417 312 35430
rect 237 35383 304 35417
rect 346 35396 422 35430
rect 338 35383 422 35396
rect 237 35358 422 35383
rect 237 35349 312 35358
rect 237 35315 304 35349
rect 346 35324 422 35358
rect 338 35315 422 35324
rect 237 35286 422 35315
rect 237 35281 312 35286
rect 237 35247 304 35281
rect 346 35252 422 35286
rect 338 35247 422 35252
rect 237 35214 422 35247
rect 237 35213 312 35214
rect 237 35179 304 35213
rect 346 35180 422 35214
rect 338 35179 422 35180
rect 237 35145 422 35179
rect 237 35111 304 35145
rect 338 35142 422 35145
rect 237 35108 312 35111
rect 346 35108 422 35142
rect 237 35077 422 35108
rect 237 35043 304 35077
rect 338 35070 422 35077
rect 237 35036 312 35043
rect 346 35036 422 35070
rect 237 35009 422 35036
rect 237 34975 304 35009
rect 338 34998 422 35009
rect 237 34964 312 34975
rect 346 34964 422 34998
rect 237 34941 422 34964
rect 237 34907 304 34941
rect 338 34926 422 34941
rect 237 34892 312 34907
rect 346 34892 422 34926
rect 237 34873 422 34892
rect 237 34839 304 34873
rect 338 34854 422 34873
rect 237 34820 312 34839
rect 346 34820 422 34854
rect 237 34805 422 34820
rect 237 34771 304 34805
rect 338 34782 422 34805
rect 237 34748 312 34771
rect 346 34748 422 34782
rect 237 34737 422 34748
rect 237 34703 304 34737
rect 338 34710 422 34737
rect 237 34676 312 34703
rect 346 34676 422 34710
rect 237 34669 422 34676
rect 237 34635 304 34669
rect 338 34638 422 34669
rect 237 34604 312 34635
rect 346 34604 422 34638
rect 237 34601 422 34604
rect 237 34567 304 34601
rect 338 34567 422 34601
rect 237 34566 422 34567
rect 237 34533 312 34566
rect 237 34499 304 34533
rect 346 34532 422 34566
rect 338 34499 422 34532
rect 237 34494 422 34499
rect 237 34465 312 34494
rect 237 34431 304 34465
rect 346 34460 422 34494
rect 338 34431 422 34460
rect 237 34422 422 34431
rect 237 34397 312 34422
rect 237 34363 304 34397
rect 346 34388 422 34422
rect 338 34363 422 34388
rect 237 34350 422 34363
rect 237 34329 312 34350
rect 237 34295 304 34329
rect 346 34316 422 34350
rect 338 34295 422 34316
rect 237 34278 422 34295
rect 237 34261 312 34278
rect 237 34227 304 34261
rect 346 34244 422 34278
rect 338 34227 422 34244
rect 237 34206 422 34227
rect 237 34193 312 34206
rect 237 34159 304 34193
rect 346 34172 422 34206
rect 338 34159 422 34172
rect 237 34134 422 34159
rect 237 34125 312 34134
rect 237 34091 304 34125
rect 346 34100 422 34134
rect 338 34091 422 34100
rect 237 34062 422 34091
rect 237 34057 312 34062
rect 237 34023 304 34057
rect 346 34028 422 34062
rect 338 34023 422 34028
rect 237 33990 422 34023
rect 237 33989 312 33990
rect 237 33955 304 33989
rect 346 33956 422 33990
rect 338 33955 422 33956
rect 237 33921 422 33955
rect 237 33887 304 33921
rect 338 33918 422 33921
rect 237 33884 312 33887
rect 346 33884 422 33918
rect 237 33853 422 33884
rect 237 33819 304 33853
rect 338 33846 422 33853
rect 237 33812 312 33819
rect 346 33812 422 33846
rect 237 33785 422 33812
rect 237 33751 304 33785
rect 338 33774 422 33785
rect 237 33740 312 33751
rect 346 33740 422 33774
rect 237 33717 422 33740
rect 237 33683 304 33717
rect 338 33702 422 33717
rect 237 33668 312 33683
rect 346 33668 422 33702
rect 237 33649 422 33668
rect 237 33615 304 33649
rect 338 33630 422 33649
rect 237 33596 312 33615
rect 346 33596 422 33630
rect 237 33581 422 33596
rect 237 33547 304 33581
rect 338 33558 422 33581
rect 237 33524 312 33547
rect 346 33524 422 33558
rect 237 33513 422 33524
rect 237 33479 304 33513
rect 338 33486 422 33513
rect 237 33452 312 33479
rect 346 33452 422 33486
rect 237 33445 422 33452
rect 237 33411 304 33445
rect 338 33414 422 33445
rect 237 33380 312 33411
rect 346 33380 422 33414
rect 237 33377 422 33380
rect 237 33343 304 33377
rect 338 33343 422 33377
rect 237 33342 422 33343
rect 237 33309 312 33342
rect 237 33275 304 33309
rect 346 33308 422 33342
rect 338 33275 422 33308
rect 237 33270 422 33275
rect 237 33241 312 33270
rect 237 33207 304 33241
rect 346 33236 422 33270
rect 338 33207 422 33236
rect 237 33198 422 33207
rect 237 33173 312 33198
rect 237 33139 304 33173
rect 346 33164 422 33198
rect 338 33139 422 33164
rect 237 33126 422 33139
rect 237 33105 312 33126
rect 237 33071 304 33105
rect 346 33092 422 33126
rect 338 33071 422 33092
rect 237 33054 422 33071
rect 237 33037 312 33054
rect 237 33003 304 33037
rect 346 33020 422 33054
rect 338 33003 422 33020
rect 237 32982 422 33003
rect 237 32969 312 32982
rect 237 32935 304 32969
rect 346 32948 422 32982
rect 338 32935 422 32948
rect 237 32910 422 32935
rect 237 32901 312 32910
rect 237 32867 304 32901
rect 346 32876 422 32910
rect 338 32867 422 32876
rect 237 32838 422 32867
rect 237 32833 312 32838
rect 237 32799 304 32833
rect 346 32804 422 32838
rect 338 32799 422 32804
rect 237 32766 422 32799
rect 237 32765 312 32766
rect 237 32731 304 32765
rect 346 32732 422 32766
rect 338 32731 422 32732
rect 237 32697 422 32731
rect 237 32663 304 32697
rect 338 32694 422 32697
rect 237 32660 312 32663
rect 346 32660 422 32694
rect 237 32629 422 32660
rect 237 32595 304 32629
rect 338 32622 422 32629
rect 237 32588 312 32595
rect 346 32588 422 32622
rect 237 32561 422 32588
rect 237 32527 304 32561
rect 338 32550 422 32561
rect 237 32516 312 32527
rect 346 32516 422 32550
rect 237 32493 422 32516
rect 237 32459 304 32493
rect 338 32478 422 32493
rect 237 32444 312 32459
rect 346 32444 422 32478
rect 237 32425 422 32444
rect 237 32391 304 32425
rect 338 32406 422 32425
rect 237 32372 312 32391
rect 346 32372 422 32406
rect 237 32357 422 32372
rect 237 32323 304 32357
rect 338 32334 422 32357
rect 237 32300 312 32323
rect 346 32300 422 32334
rect 237 32289 422 32300
rect 237 32255 304 32289
rect 338 32262 422 32289
rect 237 32228 312 32255
rect 346 32228 422 32262
rect 237 32221 422 32228
rect 237 32187 304 32221
rect 338 32190 422 32221
rect 237 32156 312 32187
rect 346 32156 422 32190
rect 237 32153 422 32156
rect 237 32119 304 32153
rect 338 32119 422 32153
rect 237 32118 422 32119
rect 237 32085 312 32118
rect 237 32051 304 32085
rect 346 32084 422 32118
rect 338 32051 422 32084
rect 237 32046 422 32051
rect 237 32017 312 32046
rect 237 31983 304 32017
rect 346 32012 422 32046
rect 338 31983 422 32012
rect 237 31974 422 31983
rect 237 31949 312 31974
rect 237 31915 304 31949
rect 346 31940 422 31974
rect 338 31915 422 31940
rect 237 31902 422 31915
rect 237 31881 312 31902
rect 237 31847 304 31881
rect 346 31868 422 31902
rect 338 31847 422 31868
rect 237 31830 422 31847
rect 237 31813 312 31830
rect 237 31779 304 31813
rect 346 31796 422 31830
rect 338 31779 422 31796
rect 237 31758 422 31779
rect 237 31745 312 31758
rect 237 31711 304 31745
rect 346 31724 422 31758
rect 338 31711 422 31724
rect 237 31686 422 31711
rect 237 31677 312 31686
rect 237 31643 304 31677
rect 346 31652 422 31686
rect 338 31643 422 31652
rect 237 31614 422 31643
rect 237 31609 312 31614
rect 237 31575 304 31609
rect 346 31580 422 31614
rect 338 31575 422 31580
rect 237 31542 422 31575
rect 237 31541 312 31542
rect 237 31507 304 31541
rect 346 31508 422 31542
rect 338 31507 422 31508
rect 237 31473 422 31507
rect 237 31439 304 31473
rect 338 31470 422 31473
rect 237 31436 312 31439
rect 346 31436 422 31470
rect 237 31405 422 31436
rect 237 31371 304 31405
rect 338 31398 422 31405
rect 237 31364 312 31371
rect 346 31364 422 31398
rect 237 31337 422 31364
rect 237 31303 304 31337
rect 338 31326 422 31337
rect 237 31292 312 31303
rect 346 31292 422 31326
rect 237 31269 422 31292
rect 237 31235 304 31269
rect 338 31254 422 31269
rect 237 31220 312 31235
rect 346 31220 422 31254
rect 237 31201 422 31220
rect 237 31167 304 31201
rect 338 31182 422 31201
rect 237 31148 312 31167
rect 346 31148 422 31182
rect 237 31133 422 31148
rect 237 31099 304 31133
rect 338 31110 422 31133
rect 237 31076 312 31099
rect 346 31076 422 31110
rect 237 31065 422 31076
rect 237 31031 304 31065
rect 338 31038 422 31065
rect 237 31004 312 31031
rect 346 31004 422 31038
rect 237 30997 422 31004
rect 237 30963 304 30997
rect 338 30966 422 30997
rect 237 30932 312 30963
rect 346 30932 422 30966
rect 237 30929 422 30932
rect 237 30895 304 30929
rect 338 30895 422 30929
rect 237 30894 422 30895
rect 237 30861 312 30894
rect 237 30827 304 30861
rect 346 30860 422 30894
rect 338 30827 422 30860
rect 237 30822 422 30827
rect 237 30793 312 30822
rect 237 30759 304 30793
rect 346 30788 422 30822
rect 338 30759 422 30788
rect 237 30750 422 30759
rect 237 30725 312 30750
rect 237 30691 304 30725
rect 346 30716 422 30750
rect 338 30691 422 30716
rect 237 30678 422 30691
rect 237 30657 312 30678
rect 237 30623 304 30657
rect 346 30644 422 30678
rect 338 30623 422 30644
rect 237 30606 422 30623
rect 237 30589 312 30606
rect 237 30555 304 30589
rect 346 30572 422 30606
rect 338 30555 422 30572
rect 237 30534 422 30555
rect 237 30521 312 30534
rect 237 30487 304 30521
rect 346 30500 422 30534
rect 338 30487 422 30500
rect 237 30462 422 30487
rect 237 30453 312 30462
rect 237 30419 304 30453
rect 346 30428 422 30462
rect 338 30419 422 30428
rect 237 30390 422 30419
rect 237 30385 312 30390
rect 237 30351 304 30385
rect 346 30356 422 30390
rect 338 30351 422 30356
rect 237 30318 422 30351
rect 237 30317 312 30318
rect 237 30283 304 30317
rect 346 30284 422 30318
rect 338 30283 422 30284
rect 237 30249 422 30283
rect 237 30215 304 30249
rect 338 30246 422 30249
rect 237 30212 312 30215
rect 346 30212 422 30246
rect 237 30181 422 30212
rect 237 30147 304 30181
rect 338 30174 422 30181
rect 237 30140 312 30147
rect 346 30140 422 30174
rect 237 30113 422 30140
rect 237 30079 304 30113
rect 338 30102 422 30113
rect 237 30068 312 30079
rect 346 30068 422 30102
rect 237 30045 422 30068
rect 237 30011 304 30045
rect 338 30030 422 30045
rect 237 29996 312 30011
rect 346 29996 422 30030
rect 237 29977 422 29996
rect 237 29943 304 29977
rect 338 29958 422 29977
rect 237 29924 312 29943
rect 346 29924 422 29958
rect 237 29909 422 29924
rect 237 29875 304 29909
rect 338 29886 422 29909
rect 237 29852 312 29875
rect 346 29852 422 29886
rect 237 29841 422 29852
rect 237 29807 304 29841
rect 338 29814 422 29841
rect 237 29780 312 29807
rect 346 29780 422 29814
rect 237 29773 422 29780
rect 237 29739 304 29773
rect 338 29742 422 29773
rect 237 29708 312 29739
rect 346 29708 422 29742
rect 237 29705 422 29708
rect 237 29671 304 29705
rect 338 29671 422 29705
rect 237 29670 422 29671
rect 237 29637 312 29670
rect 237 29603 304 29637
rect 346 29636 422 29670
rect 338 29603 422 29636
rect 237 29598 422 29603
rect 237 29569 312 29598
rect 237 29535 304 29569
rect 346 29564 422 29598
rect 338 29535 422 29564
rect 237 29526 422 29535
rect 237 29501 312 29526
rect 237 29467 304 29501
rect 346 29492 422 29526
rect 338 29467 422 29492
rect 237 29454 422 29467
rect 237 29433 312 29454
rect 237 29399 304 29433
rect 346 29420 422 29454
rect 338 29399 422 29420
rect 237 29382 422 29399
rect 237 29365 312 29382
rect 237 29331 304 29365
rect 346 29348 422 29382
rect 338 29331 422 29348
rect 237 29310 422 29331
rect 237 29297 312 29310
rect 237 29263 304 29297
rect 346 29276 422 29310
rect 338 29263 422 29276
rect 237 29238 422 29263
rect 237 29229 312 29238
rect 237 29195 304 29229
rect 346 29204 422 29238
rect 338 29195 422 29204
rect 237 29166 422 29195
rect 237 29161 312 29166
rect 237 29127 304 29161
rect 346 29132 422 29166
rect 338 29127 422 29132
rect 237 29094 422 29127
rect 237 29093 312 29094
rect 237 29059 304 29093
rect 346 29060 422 29094
rect 338 29059 422 29060
rect 237 29025 422 29059
rect 237 28991 304 29025
rect 338 29022 422 29025
rect 237 28988 312 28991
rect 346 28988 422 29022
rect 237 28957 422 28988
rect 237 28923 304 28957
rect 338 28950 422 28957
rect 237 28916 312 28923
rect 346 28916 422 28950
rect 237 28889 422 28916
rect 237 28855 304 28889
rect 338 28878 422 28889
rect 237 28844 312 28855
rect 346 28844 422 28878
rect 237 28821 422 28844
rect 237 28787 304 28821
rect 338 28806 422 28821
rect 237 28772 312 28787
rect 346 28772 422 28806
rect 237 28753 422 28772
rect 237 28719 304 28753
rect 338 28734 422 28753
rect 237 28700 312 28719
rect 346 28700 422 28734
rect 237 28685 422 28700
rect 237 28651 304 28685
rect 338 28662 422 28685
rect 237 28628 312 28651
rect 346 28628 422 28662
rect 237 28617 422 28628
rect 237 28583 304 28617
rect 338 28590 422 28617
rect 237 28556 312 28583
rect 346 28556 422 28590
rect 237 28549 422 28556
rect 237 28515 304 28549
rect 338 28518 422 28549
rect 237 28484 312 28515
rect 346 28484 422 28518
rect 237 28481 422 28484
rect 237 28447 304 28481
rect 338 28447 422 28481
rect 237 28446 422 28447
rect 237 28413 312 28446
rect 237 28379 304 28413
rect 346 28412 422 28446
rect 338 28379 422 28412
rect 237 28374 422 28379
rect 237 28345 312 28374
rect 237 28311 304 28345
rect 346 28340 422 28374
rect 338 28311 422 28340
rect 237 28302 422 28311
rect 237 28277 312 28302
rect 237 28243 304 28277
rect 346 28268 422 28302
rect 338 28243 422 28268
rect 237 28230 422 28243
rect 237 28209 312 28230
rect 237 28175 304 28209
rect 346 28196 422 28230
rect 338 28175 422 28196
rect 237 28158 422 28175
rect 237 28141 312 28158
rect 237 28107 304 28141
rect 346 28124 422 28158
rect 338 28107 422 28124
rect 237 28086 422 28107
rect 237 28073 312 28086
rect 237 28039 304 28073
rect 346 28052 422 28086
rect 338 28039 422 28052
rect 237 28014 422 28039
rect 237 28005 312 28014
rect 237 27971 304 28005
rect 346 27980 422 28014
rect 338 27971 422 27980
rect 237 27942 422 27971
rect 237 27937 312 27942
rect 237 27903 304 27937
rect 346 27908 422 27942
rect 338 27903 422 27908
rect 237 27870 422 27903
rect 237 27869 312 27870
rect 237 27835 304 27869
rect 346 27836 422 27870
rect 338 27835 422 27836
rect 237 27801 422 27835
rect 237 27767 304 27801
rect 338 27798 422 27801
rect 237 27764 312 27767
rect 346 27764 422 27798
rect 237 27733 422 27764
rect 237 27699 304 27733
rect 338 27726 422 27733
rect 237 27692 312 27699
rect 346 27692 422 27726
rect 237 27665 422 27692
rect 237 27631 304 27665
rect 338 27654 422 27665
rect 237 27620 312 27631
rect 346 27620 422 27654
rect 237 27597 422 27620
rect 237 27563 304 27597
rect 338 27582 422 27597
rect 237 27548 312 27563
rect 346 27548 422 27582
rect 237 27529 422 27548
rect 237 27495 304 27529
rect 338 27510 422 27529
rect 237 27476 312 27495
rect 346 27476 422 27510
rect 237 27461 422 27476
rect 237 27427 304 27461
rect 338 27438 422 27461
rect 237 27404 312 27427
rect 346 27404 422 27438
rect 237 27393 422 27404
rect 237 27359 304 27393
rect 338 27366 422 27393
rect 237 27332 312 27359
rect 346 27332 422 27366
rect 237 27325 422 27332
rect 237 27291 304 27325
rect 338 27294 422 27325
rect 237 27260 312 27291
rect 346 27260 422 27294
rect 237 27257 422 27260
rect 237 27223 304 27257
rect 338 27223 422 27257
rect 237 27222 422 27223
rect 237 27189 312 27222
rect 237 27155 304 27189
rect 346 27188 422 27222
rect 338 27155 422 27188
rect 237 27150 422 27155
rect 237 27121 312 27150
rect 237 27087 304 27121
rect 346 27116 422 27150
rect 338 27087 422 27116
rect 237 27078 422 27087
rect 237 27053 312 27078
rect 237 27019 304 27053
rect 346 27044 422 27078
rect 338 27019 422 27044
rect 237 27006 422 27019
rect 237 26985 312 27006
rect 237 26951 304 26985
rect 346 26972 422 27006
rect 338 26951 422 26972
rect 237 26934 422 26951
rect 237 26917 312 26934
rect 237 26883 304 26917
rect 346 26900 422 26934
rect 338 26883 422 26900
rect 237 26862 422 26883
rect 237 26849 312 26862
rect 237 26815 304 26849
rect 346 26828 422 26862
rect 338 26815 422 26828
rect 237 26790 422 26815
rect 237 26781 312 26790
rect 237 26747 304 26781
rect 346 26756 422 26790
rect 338 26747 422 26756
rect 237 26718 422 26747
rect 237 26713 312 26718
rect 237 26679 304 26713
rect 346 26684 422 26718
rect 338 26679 422 26684
rect 237 26646 422 26679
rect 237 26645 312 26646
rect 237 26611 304 26645
rect 346 26612 422 26646
rect 338 26611 422 26612
rect 237 26577 422 26611
rect 237 26543 304 26577
rect 338 26574 422 26577
rect 237 26540 312 26543
rect 346 26540 422 26574
rect 237 26509 422 26540
rect 237 26475 304 26509
rect 338 26502 422 26509
rect 237 26468 312 26475
rect 346 26468 422 26502
rect 237 26441 422 26468
rect 237 26407 304 26441
rect 338 26430 422 26441
rect 237 26396 312 26407
rect 346 26396 422 26430
rect 237 26373 422 26396
rect 237 26339 304 26373
rect 338 26358 422 26373
rect 237 26324 312 26339
rect 346 26324 422 26358
rect 237 26305 422 26324
rect 237 26271 304 26305
rect 338 26286 422 26305
rect 237 26252 312 26271
rect 346 26252 422 26286
rect 237 26237 422 26252
rect 237 26203 304 26237
rect 338 26214 422 26237
rect 237 26180 312 26203
rect 346 26180 422 26214
rect 237 26169 422 26180
rect 237 26135 304 26169
rect 338 26142 422 26169
rect 237 26108 312 26135
rect 346 26108 422 26142
rect 237 26101 422 26108
rect 237 26067 304 26101
rect 338 26070 422 26101
rect 237 26036 312 26067
rect 346 26036 422 26070
rect 237 26033 422 26036
rect 237 25999 304 26033
rect 338 25999 422 26033
rect 237 25998 422 25999
rect 237 25965 312 25998
rect 237 25931 304 25965
rect 346 25964 422 25998
rect 338 25931 422 25964
rect 237 25926 422 25931
rect 237 25897 312 25926
rect 237 25863 304 25897
rect 346 25892 422 25926
rect 338 25863 422 25892
rect 237 25854 422 25863
rect 237 25829 312 25854
rect 237 25795 304 25829
rect 346 25820 422 25854
rect 338 25795 422 25820
rect 237 25782 422 25795
rect 237 25761 312 25782
rect 237 25727 304 25761
rect 346 25748 422 25782
rect 338 25727 422 25748
rect 237 25710 422 25727
rect 237 25693 312 25710
rect 237 25659 304 25693
rect 346 25676 422 25710
rect 338 25659 422 25676
rect 237 25638 422 25659
rect 237 25625 312 25638
rect 237 25591 304 25625
rect 346 25604 422 25638
rect 338 25591 422 25604
rect 237 25566 422 25591
rect 237 25557 312 25566
rect 237 25523 304 25557
rect 346 25532 422 25566
rect 338 25523 422 25532
rect 237 25494 422 25523
rect 237 25489 312 25494
rect 237 25455 304 25489
rect 346 25460 422 25494
rect 338 25455 422 25460
rect 237 25422 422 25455
rect 237 25421 312 25422
rect 237 25387 304 25421
rect 346 25388 422 25422
rect 338 25387 422 25388
rect 237 25353 422 25387
rect 237 25319 304 25353
rect 338 25350 422 25353
rect 237 25316 312 25319
rect 346 25316 422 25350
rect 237 25285 422 25316
rect 237 25251 304 25285
rect 338 25278 422 25285
rect 237 25244 312 25251
rect 346 25244 422 25278
rect 237 25217 422 25244
rect 237 25183 304 25217
rect 338 25206 422 25217
rect 237 25172 312 25183
rect 346 25172 422 25206
rect 237 25149 422 25172
rect 237 25115 304 25149
rect 338 25134 422 25149
rect 237 25100 312 25115
rect 346 25100 422 25134
rect 237 25081 422 25100
rect 237 25047 304 25081
rect 338 25062 422 25081
rect 237 25028 312 25047
rect 346 25028 422 25062
rect 237 25013 422 25028
rect 237 24979 304 25013
rect 338 24990 422 25013
rect 237 24956 312 24979
rect 346 24956 422 24990
rect 237 24945 422 24956
rect 237 24911 304 24945
rect 338 24918 422 24945
rect 237 24884 312 24911
rect 346 24884 422 24918
rect 237 24877 422 24884
rect 237 24843 304 24877
rect 338 24846 422 24877
rect 237 24812 312 24843
rect 346 24812 422 24846
rect 237 24809 422 24812
rect 237 24775 304 24809
rect 338 24775 422 24809
rect 237 24774 422 24775
rect 237 24741 312 24774
rect 237 24707 304 24741
rect 346 24740 422 24774
rect 338 24707 422 24740
rect 237 24702 422 24707
rect 237 24673 312 24702
rect 237 24639 304 24673
rect 346 24668 422 24702
rect 338 24639 422 24668
rect 237 24630 422 24639
rect 237 24605 312 24630
rect 237 24571 304 24605
rect 346 24596 422 24630
rect 338 24571 422 24596
rect 237 24558 422 24571
rect 237 24537 312 24558
rect 237 24503 304 24537
rect 346 24524 422 24558
rect 338 24503 422 24524
rect 237 24486 422 24503
rect 237 24469 312 24486
rect 237 24435 304 24469
rect 346 24452 422 24486
rect 338 24435 422 24452
rect 237 24414 422 24435
rect 237 24401 312 24414
rect 237 24367 304 24401
rect 346 24380 422 24414
rect 338 24367 422 24380
rect 237 24342 422 24367
rect 237 24333 312 24342
rect 237 24299 304 24333
rect 346 24308 422 24342
rect 338 24299 422 24308
rect 237 24270 422 24299
rect 237 24265 312 24270
rect 237 24231 304 24265
rect 346 24236 422 24270
rect 338 24231 422 24236
rect 237 24198 422 24231
rect 237 24197 312 24198
rect 237 24163 304 24197
rect 346 24164 422 24198
rect 338 24163 422 24164
rect 237 24129 422 24163
rect 237 24095 304 24129
rect 338 24126 422 24129
rect 237 24092 312 24095
rect 346 24092 422 24126
rect 237 24061 422 24092
rect 237 24027 304 24061
rect 338 24054 422 24061
rect 237 24020 312 24027
rect 346 24020 422 24054
rect 237 23993 422 24020
rect 237 23959 304 23993
rect 338 23982 422 23993
rect 237 23948 312 23959
rect 346 23948 422 23982
rect 237 23925 422 23948
rect 237 23891 304 23925
rect 338 23910 422 23925
rect 237 23876 312 23891
rect 346 23876 422 23910
rect 237 23857 422 23876
rect 237 23823 304 23857
rect 338 23838 422 23857
rect 237 23804 312 23823
rect 346 23804 422 23838
rect 237 23789 422 23804
rect 237 23755 304 23789
rect 338 23766 422 23789
rect 237 23732 312 23755
rect 346 23732 422 23766
rect 237 23721 422 23732
rect 237 23687 304 23721
rect 338 23694 422 23721
rect 237 23660 312 23687
rect 346 23660 422 23694
rect 237 23653 422 23660
rect 237 23619 304 23653
rect 338 23622 422 23653
rect 237 23588 312 23619
rect 346 23588 422 23622
rect 237 23585 422 23588
rect 237 23551 304 23585
rect 338 23551 422 23585
rect 237 23550 422 23551
rect 237 23517 312 23550
rect 237 23483 304 23517
rect 346 23516 422 23550
rect 338 23483 422 23516
rect 237 23478 422 23483
rect 237 23449 312 23478
rect 237 23415 304 23449
rect 346 23444 422 23478
rect 338 23415 422 23444
rect 237 23406 422 23415
rect 237 23381 312 23406
rect 237 23347 304 23381
rect 346 23372 422 23406
rect 338 23347 422 23372
rect 237 23334 422 23347
rect 237 23313 312 23334
rect 237 23279 304 23313
rect 346 23300 422 23334
rect 338 23279 422 23300
rect 237 23262 422 23279
rect 237 23245 312 23262
rect 237 23211 304 23245
rect 346 23228 422 23262
rect 338 23211 422 23228
rect 237 23190 422 23211
rect 237 23177 312 23190
rect 237 23143 304 23177
rect 346 23156 422 23190
rect 338 23143 422 23156
rect 237 23118 422 23143
rect 237 23109 312 23118
rect 237 23075 304 23109
rect 346 23084 422 23118
rect 338 23075 422 23084
rect 237 23046 422 23075
rect 237 23041 312 23046
rect 237 23007 304 23041
rect 346 23012 422 23046
rect 338 23007 422 23012
rect 237 22974 422 23007
rect 237 22973 312 22974
rect 237 22939 304 22973
rect 346 22940 422 22974
rect 338 22939 422 22940
rect 237 22905 422 22939
rect 237 22871 304 22905
rect 338 22902 422 22905
rect 237 22868 312 22871
rect 346 22868 422 22902
rect 237 22837 422 22868
rect 237 22803 304 22837
rect 338 22830 422 22837
rect 237 22796 312 22803
rect 346 22796 422 22830
rect 237 22769 422 22796
rect 237 22735 304 22769
rect 338 22758 422 22769
rect 237 22724 312 22735
rect 346 22724 422 22758
rect 237 22701 422 22724
rect 237 22667 304 22701
rect 338 22686 422 22701
rect 237 22652 312 22667
rect 346 22652 422 22686
rect 237 22633 422 22652
rect 237 22599 304 22633
rect 338 22614 422 22633
rect 237 22580 312 22599
rect 346 22580 422 22614
rect 237 22565 422 22580
rect 237 22531 304 22565
rect 338 22542 422 22565
rect 237 22508 312 22531
rect 346 22508 422 22542
rect 237 22497 422 22508
rect 237 22463 304 22497
rect 338 22470 422 22497
rect 237 22436 312 22463
rect 346 22436 422 22470
rect 237 22429 422 22436
rect 237 22395 304 22429
rect 338 22398 422 22429
rect 237 22364 312 22395
rect 346 22364 422 22398
rect 237 22361 422 22364
rect 237 22327 304 22361
rect 338 22327 422 22361
rect 237 22326 422 22327
rect 237 22293 312 22326
rect 237 22259 304 22293
rect 346 22292 422 22326
rect 338 22259 422 22292
rect 237 22254 422 22259
rect 237 22225 312 22254
rect 237 22191 304 22225
rect 346 22220 422 22254
rect 338 22191 422 22220
rect 237 22182 422 22191
rect 237 22157 312 22182
rect 237 22123 304 22157
rect 346 22148 422 22182
rect 338 22123 422 22148
rect 237 22110 422 22123
rect 237 22089 312 22110
rect 237 22055 304 22089
rect 346 22076 422 22110
rect 338 22055 422 22076
rect 237 22038 422 22055
rect 237 22021 312 22038
rect 237 21987 304 22021
rect 346 22004 422 22038
rect 338 21987 422 22004
rect 237 21966 422 21987
rect 237 21953 312 21966
rect 237 21919 304 21953
rect 346 21932 422 21966
rect 338 21919 422 21932
rect 237 21894 422 21919
rect 237 21885 312 21894
rect 237 21851 304 21885
rect 346 21860 422 21894
rect 338 21851 422 21860
rect 237 21822 422 21851
rect 237 21817 312 21822
rect 237 21783 304 21817
rect 346 21788 422 21822
rect 338 21783 422 21788
rect 237 21750 422 21783
rect 237 21749 312 21750
rect 237 21715 304 21749
rect 346 21716 422 21750
rect 338 21715 422 21716
rect 237 21681 422 21715
rect 237 21647 304 21681
rect 338 21678 422 21681
rect 237 21644 312 21647
rect 346 21644 422 21678
rect 237 21613 422 21644
rect 237 21579 304 21613
rect 338 21606 422 21613
rect 237 21572 312 21579
rect 346 21572 422 21606
rect 237 21545 422 21572
rect 237 21511 304 21545
rect 338 21534 422 21545
rect 237 21500 312 21511
rect 346 21500 422 21534
rect 237 21477 422 21500
rect 237 21443 304 21477
rect 338 21462 422 21477
rect 237 21428 312 21443
rect 346 21428 422 21462
rect 237 21409 422 21428
rect 237 21375 304 21409
rect 338 21390 422 21409
rect 237 21356 312 21375
rect 346 21356 422 21390
rect 237 21341 422 21356
rect 237 21307 304 21341
rect 338 21318 422 21341
rect 237 21284 312 21307
rect 346 21284 422 21318
rect 237 21273 422 21284
rect 237 21239 304 21273
rect 338 21246 422 21273
rect 237 21212 312 21239
rect 346 21212 422 21246
rect 237 21205 422 21212
rect 237 21171 304 21205
rect 338 21174 422 21205
rect 237 21140 312 21171
rect 346 21140 422 21174
rect 237 21137 422 21140
rect 237 21103 304 21137
rect 338 21103 422 21137
rect 237 21102 422 21103
rect 237 21069 312 21102
rect 237 21035 304 21069
rect 346 21068 422 21102
rect 338 21035 422 21068
rect 237 21030 422 21035
rect 237 21001 312 21030
rect 237 20967 304 21001
rect 346 20996 422 21030
rect 338 20967 422 20996
rect 237 20958 422 20967
rect 237 20933 312 20958
rect 237 20899 304 20933
rect 346 20924 422 20958
rect 338 20899 422 20924
rect 237 20886 422 20899
rect 237 20865 312 20886
rect 237 20831 304 20865
rect 346 20852 422 20886
rect 338 20831 422 20852
rect 237 20814 422 20831
rect 237 20797 312 20814
rect 237 20763 304 20797
rect 346 20780 422 20814
rect 338 20763 422 20780
rect 237 20742 422 20763
rect 237 20729 312 20742
rect 237 20695 304 20729
rect 346 20708 422 20742
rect 338 20695 422 20708
rect 237 20670 422 20695
rect 237 20661 312 20670
rect 237 20627 304 20661
rect 346 20636 422 20670
rect 338 20627 422 20636
rect 237 20598 422 20627
rect 237 20593 312 20598
rect 237 20559 304 20593
rect 346 20564 422 20598
rect 338 20559 422 20564
rect 237 20526 422 20559
rect 237 20525 312 20526
rect 237 20491 304 20525
rect 346 20492 422 20526
rect 338 20491 422 20492
rect 237 20457 422 20491
rect 237 20423 304 20457
rect 338 20454 422 20457
rect 237 20420 312 20423
rect 346 20420 422 20454
rect 237 20389 422 20420
rect 237 20355 304 20389
rect 338 20382 422 20389
rect 237 20348 312 20355
rect 346 20348 422 20382
rect 237 20321 422 20348
rect 237 20287 304 20321
rect 338 20310 422 20321
rect 237 20276 312 20287
rect 346 20276 422 20310
rect 237 20253 422 20276
rect 237 20219 304 20253
rect 338 20238 422 20253
rect 237 20204 312 20219
rect 346 20204 422 20238
rect 237 20185 422 20204
rect 237 20151 304 20185
rect 338 20166 422 20185
rect 237 20132 312 20151
rect 346 20132 422 20166
rect 237 20117 422 20132
rect 237 20083 304 20117
rect 338 20094 422 20117
rect 237 20060 312 20083
rect 346 20060 422 20094
rect 237 20049 422 20060
rect 237 20015 304 20049
rect 338 20022 422 20049
rect 237 19988 312 20015
rect 346 19988 422 20022
rect 237 19981 422 19988
rect 237 19947 304 19981
rect 338 19950 422 19981
rect 237 19916 312 19947
rect 346 19916 422 19950
rect 237 19913 422 19916
rect 237 19879 304 19913
rect 338 19879 422 19913
rect 237 19878 422 19879
rect 237 19845 312 19878
rect 237 19811 304 19845
rect 346 19844 422 19878
rect 338 19811 422 19844
rect 237 19806 422 19811
rect 237 19777 312 19806
rect 237 19743 304 19777
rect 346 19772 422 19806
rect 338 19743 422 19772
rect 237 19734 422 19743
rect 237 19709 312 19734
rect 237 19675 304 19709
rect 346 19700 422 19734
rect 338 19675 422 19700
rect 237 19662 422 19675
rect 237 19641 312 19662
rect 237 19607 304 19641
rect 346 19628 422 19662
rect 338 19607 422 19628
rect 237 19590 422 19607
rect 237 19573 312 19590
rect 237 19539 304 19573
rect 346 19556 422 19590
rect 338 19539 422 19556
rect 237 19518 422 19539
rect 237 19505 312 19518
rect 237 19471 304 19505
rect 346 19484 422 19518
rect 338 19471 422 19484
rect 237 19446 422 19471
rect 237 19437 312 19446
rect 237 19403 304 19437
rect 346 19412 422 19446
rect 338 19403 422 19412
rect 237 19374 422 19403
rect 237 19369 312 19374
rect 237 19335 304 19369
rect 346 19340 422 19374
rect 338 19335 422 19340
rect 237 19302 422 19335
rect 237 19301 312 19302
rect 237 19267 304 19301
rect 346 19268 422 19302
rect 338 19267 422 19268
rect 237 19233 422 19267
rect 237 19199 304 19233
rect 338 19230 422 19233
rect 237 19196 312 19199
rect 346 19196 422 19230
rect 237 19165 422 19196
rect 237 19131 304 19165
rect 338 19158 422 19165
rect 237 19124 312 19131
rect 346 19124 422 19158
rect 237 19097 422 19124
rect 237 19063 304 19097
rect 338 19086 422 19097
rect 237 19052 312 19063
rect 346 19052 422 19086
rect 237 19029 422 19052
rect 237 18995 304 19029
rect 338 19014 422 19029
rect 237 18980 312 18995
rect 346 18980 422 19014
rect 237 18961 422 18980
rect 237 18927 304 18961
rect 338 18942 422 18961
rect 237 18908 312 18927
rect 346 18908 422 18942
rect 237 18893 422 18908
rect 237 18859 304 18893
rect 338 18870 422 18893
rect 237 18836 312 18859
rect 346 18836 422 18870
rect 237 18825 422 18836
rect 237 18791 304 18825
rect 338 18798 422 18825
rect 237 18764 312 18791
rect 346 18764 422 18798
rect 237 18757 422 18764
rect 237 18723 304 18757
rect 338 18726 422 18757
rect 237 18692 312 18723
rect 346 18692 422 18726
rect 237 18689 422 18692
rect 237 18655 304 18689
rect 338 18655 422 18689
rect 237 18654 422 18655
rect 237 18621 312 18654
rect 237 18587 304 18621
rect 346 18620 422 18654
rect 338 18587 422 18620
rect 237 18582 422 18587
rect 237 18553 312 18582
rect 237 18519 304 18553
rect 346 18548 422 18582
rect 338 18519 422 18548
rect 237 18510 422 18519
rect 237 18485 312 18510
rect 237 18451 304 18485
rect 346 18476 422 18510
rect 338 18451 422 18476
rect 237 18438 422 18451
rect 237 18417 312 18438
rect 237 18383 304 18417
rect 346 18404 422 18438
rect 338 18383 422 18404
rect 237 18366 422 18383
rect 237 18349 312 18366
rect 237 18315 304 18349
rect 346 18332 422 18366
rect 338 18315 422 18332
rect 237 18294 422 18315
rect 237 18281 312 18294
rect 237 18247 304 18281
rect 346 18260 422 18294
rect 338 18247 422 18260
rect 237 18222 422 18247
rect 237 18213 312 18222
rect 237 18179 304 18213
rect 346 18188 422 18222
rect 338 18179 422 18188
rect 237 18150 422 18179
rect 237 18145 312 18150
rect 237 18111 304 18145
rect 346 18116 422 18150
rect 338 18111 422 18116
rect 237 18078 422 18111
rect 237 18077 312 18078
rect 237 18043 304 18077
rect 346 18044 422 18078
rect 338 18043 422 18044
rect 237 18009 422 18043
rect 237 17975 304 18009
rect 338 18006 422 18009
rect 237 17972 312 17975
rect 346 17972 422 18006
rect 237 17941 422 17972
rect 237 17907 304 17941
rect 338 17934 422 17941
rect 237 17900 312 17907
rect 346 17900 422 17934
rect 237 17873 422 17900
rect 237 17839 304 17873
rect 338 17862 422 17873
rect 237 17828 312 17839
rect 346 17828 422 17862
rect 237 17805 422 17828
rect 237 17771 304 17805
rect 338 17790 422 17805
rect 237 17756 312 17771
rect 346 17756 422 17790
rect 237 17737 422 17756
rect 237 17703 304 17737
rect 338 17718 422 17737
rect 237 17684 312 17703
rect 346 17684 422 17718
rect 237 17669 422 17684
rect 237 17635 304 17669
rect 338 17646 422 17669
rect 237 17612 312 17635
rect 346 17612 422 17646
rect 237 17601 422 17612
rect 237 17567 304 17601
rect 338 17574 422 17601
rect 237 17540 312 17567
rect 346 17540 422 17574
rect 237 17533 422 17540
rect 237 17499 304 17533
rect 338 17502 422 17533
rect 237 17468 312 17499
rect 346 17468 422 17502
rect 237 17465 422 17468
rect 237 17431 304 17465
rect 338 17431 422 17465
rect 237 17430 422 17431
rect 237 17397 312 17430
rect 237 17363 304 17397
rect 346 17396 422 17430
rect 338 17363 422 17396
rect 237 17358 422 17363
rect 237 17329 312 17358
rect 237 17295 304 17329
rect 346 17324 422 17358
rect 338 17295 422 17324
rect 237 17286 422 17295
rect 237 17261 312 17286
rect 237 17227 304 17261
rect 346 17252 422 17286
rect 338 17227 422 17252
rect 237 17214 422 17227
rect 237 17193 312 17214
rect 237 17159 304 17193
rect 346 17180 422 17214
rect 338 17159 422 17180
rect 237 17142 422 17159
rect 237 17125 312 17142
rect 237 17091 304 17125
rect 346 17108 422 17142
rect 338 17091 422 17108
rect 237 17070 422 17091
rect 237 17057 312 17070
rect 237 17023 304 17057
rect 346 17036 422 17070
rect 338 17023 422 17036
rect 237 16998 422 17023
rect 237 16989 312 16998
rect 237 16955 304 16989
rect 346 16964 422 16998
rect 338 16955 422 16964
rect 237 16926 422 16955
rect 237 16921 312 16926
rect 237 16887 304 16921
rect 346 16892 422 16926
rect 338 16887 422 16892
rect 237 16854 422 16887
rect 237 16853 312 16854
rect 237 16819 304 16853
rect 346 16820 422 16854
rect 338 16819 422 16820
rect 237 16785 422 16819
rect 237 16751 304 16785
rect 338 16782 422 16785
rect 237 16748 312 16751
rect 346 16748 422 16782
rect 237 16717 422 16748
rect 237 16683 304 16717
rect 338 16710 422 16717
rect 237 16676 312 16683
rect 346 16676 422 16710
rect 237 16649 422 16676
rect 237 16615 304 16649
rect 338 16638 422 16649
rect 237 16604 312 16615
rect 346 16604 422 16638
rect 237 16581 422 16604
rect 237 16547 304 16581
rect 338 16566 422 16581
rect 237 16532 312 16547
rect 346 16532 422 16566
rect 237 16513 422 16532
rect 237 16479 304 16513
rect 338 16494 422 16513
rect 237 16460 312 16479
rect 346 16460 422 16494
rect 237 16445 422 16460
rect 237 16411 304 16445
rect 338 16422 422 16445
rect 237 16388 312 16411
rect 346 16388 422 16422
rect 237 16377 422 16388
rect 237 16343 304 16377
rect 338 16350 422 16377
rect 237 16316 312 16343
rect 346 16316 422 16350
rect 237 16309 422 16316
rect 237 16275 304 16309
rect 338 16278 422 16309
rect 237 16244 312 16275
rect 346 16244 422 16278
rect 237 16241 422 16244
rect 237 16207 304 16241
rect 338 16207 422 16241
rect 237 16206 422 16207
rect 237 16173 312 16206
rect 237 16139 304 16173
rect 346 16172 422 16206
rect 338 16139 422 16172
rect 237 16134 422 16139
rect 237 16105 312 16134
rect 237 16071 304 16105
rect 346 16100 422 16134
rect 338 16071 422 16100
rect 237 16062 422 16071
rect 237 16037 312 16062
rect 237 16003 304 16037
rect 346 16028 422 16062
rect 338 16003 422 16028
rect 237 15990 422 16003
rect 237 15969 312 15990
rect 237 15935 304 15969
rect 346 15956 422 15990
rect 338 15935 422 15956
rect 237 15918 422 15935
rect 237 15901 312 15918
rect 237 15867 304 15901
rect 346 15884 422 15918
rect 338 15867 422 15884
rect 237 15846 422 15867
rect 237 15833 312 15846
rect 237 15799 304 15833
rect 346 15812 422 15846
rect 338 15799 422 15812
rect 237 15774 422 15799
rect 237 15765 312 15774
rect 237 15731 304 15765
rect 346 15740 422 15774
rect 338 15731 422 15740
rect 237 15702 422 15731
rect 237 15697 312 15702
rect 237 15663 304 15697
rect 346 15668 422 15702
rect 338 15663 422 15668
rect 237 15630 422 15663
rect 237 15629 312 15630
rect 237 15595 304 15629
rect 346 15596 422 15630
rect 338 15595 422 15596
rect 237 15561 422 15595
rect 237 15527 304 15561
rect 338 15558 422 15561
rect 237 15524 312 15527
rect 346 15524 422 15558
rect 237 15493 422 15524
rect 237 15459 304 15493
rect 338 15486 422 15493
rect 237 15452 312 15459
rect 346 15452 422 15486
rect 237 15425 422 15452
rect 237 15391 304 15425
rect 338 15414 422 15425
rect 237 15380 312 15391
rect 346 15380 422 15414
rect 237 15357 422 15380
rect 237 15323 304 15357
rect 338 15342 422 15357
rect 237 15308 312 15323
rect 346 15308 422 15342
rect 237 15289 422 15308
rect 237 15255 304 15289
rect 338 15270 422 15289
rect 237 15236 312 15255
rect 346 15236 422 15270
rect 237 15221 422 15236
rect 237 15187 304 15221
rect 338 15198 422 15221
rect 237 15164 312 15187
rect 346 15164 422 15198
rect 237 15153 422 15164
rect 237 15119 304 15153
rect 338 15126 422 15153
rect 237 15092 312 15119
rect 346 15092 422 15126
rect 237 15085 422 15092
rect 237 15051 304 15085
rect 338 15054 422 15085
rect 237 15020 312 15051
rect 346 15020 422 15054
rect 237 15017 422 15020
rect 237 14983 304 15017
rect 338 14983 422 15017
rect 237 14982 422 14983
rect 237 14949 312 14982
rect 237 14915 304 14949
rect 346 14948 422 14982
rect 338 14915 422 14948
rect 237 14910 422 14915
rect 237 14881 312 14910
rect 237 14847 304 14881
rect 346 14876 422 14910
rect 338 14847 422 14876
rect 237 14838 422 14847
rect 237 14813 312 14838
rect 237 14779 304 14813
rect 346 14804 422 14838
rect 338 14779 422 14804
rect 237 14766 422 14779
rect 237 14745 312 14766
rect 237 14711 304 14745
rect 346 14732 422 14766
rect 338 14711 422 14732
rect 595 36190 14353 36220
rect 595 36156 758 36190
rect 792 36156 826 36190
rect 860 36156 894 36190
rect 928 36156 962 36190
rect 996 36156 1030 36190
rect 1064 36156 1098 36190
rect 1132 36156 1166 36190
rect 1200 36156 1234 36190
rect 1268 36156 1302 36190
rect 1336 36156 1370 36190
rect 1404 36156 1438 36190
rect 1472 36156 1506 36190
rect 1540 36156 1574 36190
rect 1608 36156 1642 36190
rect 1676 36156 1710 36190
rect 1744 36156 1778 36190
rect 1812 36156 1846 36190
rect 1880 36156 1914 36190
rect 1948 36156 1982 36190
rect 2016 36156 2050 36190
rect 2084 36156 2118 36190
rect 2152 36156 2186 36190
rect 2220 36156 2254 36190
rect 2288 36156 2322 36190
rect 2356 36156 2390 36190
rect 2424 36156 2458 36190
rect 2492 36156 2526 36190
rect 2560 36156 2594 36190
rect 2628 36156 2662 36190
rect 2696 36156 2730 36190
rect 2764 36156 2798 36190
rect 2832 36156 2866 36190
rect 2900 36156 2934 36190
rect 2968 36156 3002 36190
rect 3036 36156 3070 36190
rect 3104 36156 3138 36190
rect 3172 36156 3206 36190
rect 3240 36156 3274 36190
rect 3308 36156 3342 36190
rect 3376 36156 3410 36190
rect 3444 36156 3478 36190
rect 3512 36156 3546 36190
rect 3580 36156 3614 36190
rect 3648 36156 3682 36190
rect 3716 36156 3750 36190
rect 3784 36156 3818 36190
rect 3852 36156 3886 36190
rect 3920 36156 3954 36190
rect 3988 36156 4022 36190
rect 4056 36156 4090 36190
rect 4124 36156 4158 36190
rect 4192 36156 4226 36190
rect 4260 36156 4294 36190
rect 4328 36156 4362 36190
rect 4396 36156 4430 36190
rect 4464 36156 4498 36190
rect 4532 36156 4566 36190
rect 4600 36156 4634 36190
rect 4668 36156 4702 36190
rect 4736 36156 4770 36190
rect 4804 36156 4838 36190
rect 4872 36156 4906 36190
rect 4940 36156 4974 36190
rect 5008 36156 5042 36190
rect 5076 36156 5110 36190
rect 5144 36156 5178 36190
rect 5212 36156 5246 36190
rect 5280 36156 5314 36190
rect 5348 36156 5382 36190
rect 5416 36156 5450 36190
rect 5484 36156 5518 36190
rect 5552 36156 5586 36190
rect 5620 36156 5654 36190
rect 5688 36156 5722 36190
rect 5756 36156 5790 36190
rect 5824 36156 5858 36190
rect 5892 36156 5926 36190
rect 5960 36156 5994 36190
rect 6028 36156 6062 36190
rect 6096 36156 6130 36190
rect 6164 36156 6198 36190
rect 6232 36156 6266 36190
rect 6300 36156 6334 36190
rect 6368 36156 6402 36190
rect 6436 36156 6470 36190
rect 6504 36156 6538 36190
rect 6572 36156 6606 36190
rect 6640 36156 6674 36190
rect 6708 36156 6742 36190
rect 6776 36156 6810 36190
rect 6844 36156 6878 36190
rect 6912 36156 6946 36190
rect 6980 36156 7014 36190
rect 7048 36156 7082 36190
rect 7116 36156 7150 36190
rect 7184 36156 7218 36190
rect 7252 36156 7286 36190
rect 7320 36156 7354 36190
rect 7388 36156 7422 36190
rect 7456 36156 7490 36190
rect 7524 36156 7558 36190
rect 7592 36156 7626 36190
rect 7660 36156 7694 36190
rect 7728 36156 7762 36190
rect 7796 36156 7830 36190
rect 7864 36156 7898 36190
rect 7932 36156 7966 36190
rect 8000 36156 8034 36190
rect 8068 36156 8102 36190
rect 8136 36156 8170 36190
rect 8204 36156 8238 36190
rect 8272 36156 8306 36190
rect 8340 36156 8374 36190
rect 8408 36156 8442 36190
rect 8476 36156 8510 36190
rect 8544 36156 8578 36190
rect 8612 36156 8646 36190
rect 8680 36156 8714 36190
rect 8748 36156 8782 36190
rect 8816 36156 8850 36190
rect 8884 36156 8918 36190
rect 8952 36156 8986 36190
rect 9020 36156 9054 36190
rect 9088 36156 9122 36190
rect 9156 36156 9190 36190
rect 9224 36156 9258 36190
rect 9292 36156 9326 36190
rect 9360 36156 9394 36190
rect 9428 36156 9462 36190
rect 9496 36156 9530 36190
rect 9564 36156 9598 36190
rect 9632 36156 9666 36190
rect 9700 36156 9734 36190
rect 9768 36156 9802 36190
rect 9836 36156 9870 36190
rect 9904 36156 9938 36190
rect 9972 36156 10006 36190
rect 10040 36156 10074 36190
rect 10108 36156 10142 36190
rect 10176 36156 10210 36190
rect 10244 36156 10278 36190
rect 10312 36156 10346 36190
rect 10380 36156 10414 36190
rect 10448 36156 10482 36190
rect 10516 36156 10550 36190
rect 10584 36156 10618 36190
rect 10652 36156 10686 36190
rect 10720 36156 10754 36190
rect 10788 36156 10822 36190
rect 10856 36156 10890 36190
rect 10924 36156 10958 36190
rect 10992 36156 11026 36190
rect 11060 36156 11094 36190
rect 11128 36156 11162 36190
rect 11196 36156 11230 36190
rect 11264 36156 11298 36190
rect 11332 36156 11366 36190
rect 11400 36156 11434 36190
rect 11468 36156 11502 36190
rect 11536 36156 11570 36190
rect 11604 36156 11638 36190
rect 11672 36156 11706 36190
rect 11740 36156 11774 36190
rect 11808 36156 11842 36190
rect 11876 36156 11910 36190
rect 11944 36156 11978 36190
rect 12012 36156 12046 36190
rect 12080 36156 12114 36190
rect 12148 36156 12182 36190
rect 12216 36156 12250 36190
rect 12284 36156 12318 36190
rect 12352 36156 12386 36190
rect 12420 36156 12454 36190
rect 12488 36156 12522 36190
rect 12556 36156 12590 36190
rect 12624 36156 12658 36190
rect 12692 36156 12726 36190
rect 12760 36156 12794 36190
rect 12828 36156 12862 36190
rect 12896 36156 12930 36190
rect 12964 36156 12998 36190
rect 13032 36156 13066 36190
rect 13100 36156 13134 36190
rect 13168 36156 13202 36190
rect 13236 36156 13270 36190
rect 13304 36156 13338 36190
rect 13372 36156 13406 36190
rect 13440 36156 13474 36190
rect 13508 36156 13542 36190
rect 13576 36156 13610 36190
rect 13644 36156 13678 36190
rect 13712 36156 13746 36190
rect 13780 36156 13814 36190
rect 13848 36156 13882 36190
rect 13916 36156 13950 36190
rect 13984 36156 14018 36190
rect 14052 36156 14086 36190
rect 14120 36156 14154 36190
rect 14188 36156 14353 36190
rect 595 36063 14353 36156
rect 595 36029 624 36063
rect 658 36029 14289 36063
rect 14323 36029 14353 36063
rect 595 36016 14353 36029
rect 595 35995 1001 36016
rect 595 35961 624 35995
rect 658 35982 1001 35995
rect 1035 35982 1073 36016
rect 1107 35982 1145 36016
rect 1179 35982 1217 36016
rect 1251 35982 1289 36016
rect 1323 35982 1361 36016
rect 1395 35982 1433 36016
rect 1467 35982 1505 36016
rect 1539 35982 1577 36016
rect 1611 35982 1649 36016
rect 1683 35982 1721 36016
rect 1755 35982 1793 36016
rect 1827 35982 1865 36016
rect 1899 35982 1937 36016
rect 1971 35982 2009 36016
rect 2043 35982 2081 36016
rect 2115 35982 2153 36016
rect 2187 35982 2225 36016
rect 2259 35982 2297 36016
rect 2331 35982 2369 36016
rect 2403 35982 2441 36016
rect 2475 35982 2513 36016
rect 2547 35982 2585 36016
rect 2619 35982 2657 36016
rect 2691 35982 2729 36016
rect 2763 35982 2801 36016
rect 2835 35982 2873 36016
rect 2907 35982 2945 36016
rect 2979 35982 3017 36016
rect 3051 35982 3089 36016
rect 3123 35982 3161 36016
rect 3195 35982 3233 36016
rect 3267 35982 3305 36016
rect 3339 35982 3377 36016
rect 3411 35982 3449 36016
rect 3483 35982 3521 36016
rect 3555 35982 3593 36016
rect 3627 35982 3665 36016
rect 3699 35982 3737 36016
rect 3771 35982 3809 36016
rect 3843 35982 3881 36016
rect 3915 35982 3953 36016
rect 3987 35982 4025 36016
rect 4059 35982 4097 36016
rect 4131 35982 4169 36016
rect 4203 35982 4241 36016
rect 4275 35982 4313 36016
rect 4347 35982 4385 36016
rect 4419 35982 4457 36016
rect 4491 35982 4529 36016
rect 4563 35982 4601 36016
rect 4635 35982 4673 36016
rect 4707 35982 4745 36016
rect 4779 35982 4817 36016
rect 4851 35982 4889 36016
rect 4923 35982 4961 36016
rect 4995 35982 5033 36016
rect 5067 35982 5105 36016
rect 5139 35982 5177 36016
rect 5211 35982 5249 36016
rect 5283 35982 5321 36016
rect 5355 35982 5393 36016
rect 5427 35982 5465 36016
rect 5499 35982 5537 36016
rect 5571 35982 5609 36016
rect 5643 35982 5681 36016
rect 5715 35982 5753 36016
rect 5787 35982 5825 36016
rect 5859 35982 5897 36016
rect 5931 35982 5969 36016
rect 6003 35982 6041 36016
rect 6075 35982 6113 36016
rect 6147 35982 6185 36016
rect 6219 35982 6257 36016
rect 6291 35982 6329 36016
rect 6363 35982 6401 36016
rect 6435 35982 6473 36016
rect 6507 35982 6545 36016
rect 6579 35982 6617 36016
rect 6651 35982 6689 36016
rect 6723 35982 6761 36016
rect 6795 35982 6833 36016
rect 6867 35982 6905 36016
rect 6939 35982 6977 36016
rect 7011 35982 7049 36016
rect 7083 35982 7121 36016
rect 7155 35982 7193 36016
rect 7227 35982 7265 36016
rect 7299 35982 7337 36016
rect 7371 35982 7409 36016
rect 7443 35982 7481 36016
rect 7515 35982 7553 36016
rect 7587 35982 7625 36016
rect 7659 35982 7697 36016
rect 7731 35982 7769 36016
rect 7803 35982 7841 36016
rect 7875 35982 7913 36016
rect 7947 35982 7985 36016
rect 8019 35982 8057 36016
rect 8091 35982 8129 36016
rect 8163 35982 8201 36016
rect 8235 35982 8273 36016
rect 8307 35982 8345 36016
rect 8379 35982 8417 36016
rect 8451 35982 8489 36016
rect 8523 35982 8561 36016
rect 8595 35982 8633 36016
rect 8667 35982 8705 36016
rect 8739 35982 8777 36016
rect 8811 35982 8849 36016
rect 8883 35982 8921 36016
rect 8955 35982 8993 36016
rect 9027 35982 9065 36016
rect 9099 35982 9137 36016
rect 9171 35982 9209 36016
rect 9243 35982 9281 36016
rect 9315 35982 9353 36016
rect 9387 35982 9425 36016
rect 9459 35982 9497 36016
rect 9531 35982 9569 36016
rect 9603 35982 9641 36016
rect 9675 35982 9713 36016
rect 9747 35982 9785 36016
rect 9819 35982 9857 36016
rect 9891 35982 9929 36016
rect 9963 35982 10001 36016
rect 10035 35982 10073 36016
rect 10107 35982 10145 36016
rect 10179 35982 10217 36016
rect 10251 35982 10289 36016
rect 10323 35982 10361 36016
rect 10395 35982 10433 36016
rect 10467 35982 10505 36016
rect 10539 35982 10577 36016
rect 10611 35982 10649 36016
rect 10683 35982 10721 36016
rect 10755 35982 10793 36016
rect 10827 35982 10865 36016
rect 10899 35982 10937 36016
rect 10971 35982 11009 36016
rect 11043 35982 11081 36016
rect 11115 35982 11153 36016
rect 11187 35982 11225 36016
rect 11259 35982 11297 36016
rect 11331 35982 11369 36016
rect 11403 35982 11441 36016
rect 11475 35982 11513 36016
rect 11547 35982 11585 36016
rect 11619 35982 11657 36016
rect 11691 35982 11729 36016
rect 11763 35982 11801 36016
rect 11835 35982 11873 36016
rect 11907 35982 11945 36016
rect 11979 35982 12017 36016
rect 12051 35982 12089 36016
rect 12123 35982 12161 36016
rect 12195 35982 12233 36016
rect 12267 35982 12305 36016
rect 12339 35982 12377 36016
rect 12411 35982 12449 36016
rect 12483 35982 12521 36016
rect 12555 35982 12593 36016
rect 12627 35982 12665 36016
rect 12699 35982 12737 36016
rect 12771 35982 12809 36016
rect 12843 35982 12881 36016
rect 12915 35982 12953 36016
rect 12987 35982 13025 36016
rect 13059 35982 13097 36016
rect 13131 35982 13169 36016
rect 13203 35982 13241 36016
rect 13275 35982 13313 36016
rect 13347 35982 13385 36016
rect 13419 35982 13457 36016
rect 13491 35982 13529 36016
rect 13563 35982 13601 36016
rect 13635 35982 13673 36016
rect 13707 35982 13745 36016
rect 13779 35982 13817 36016
rect 13851 35982 13889 36016
rect 13923 35982 13961 36016
rect 13995 35995 14353 36016
rect 13995 35982 14289 35995
rect 658 35961 14289 35982
rect 14323 35961 14353 35995
rect 595 35927 14353 35961
rect 595 35893 624 35927
rect 658 35913 14289 35927
rect 658 35893 799 35913
rect 595 35879 799 35893
rect 833 35893 14289 35913
rect 14323 35893 14353 35927
rect 833 35879 14353 35893
rect 595 35859 14353 35879
rect 595 35825 624 35859
rect 658 35841 14289 35859
rect 658 35825 799 35841
rect 595 35807 799 35825
rect 833 35834 14289 35841
rect 833 35807 14114 35834
rect 595 35800 14114 35807
rect 14148 35825 14289 35834
rect 14323 35825 14353 35859
rect 14148 35800 14353 35825
rect 595 35791 14353 35800
rect 595 35757 624 35791
rect 658 35769 14289 35791
rect 658 35757 799 35769
rect 595 35735 799 35757
rect 833 35762 14289 35769
rect 833 35735 14114 35762
rect 595 35728 14114 35735
rect 14148 35757 14289 35762
rect 14323 35757 14353 35791
rect 14148 35728 14353 35757
rect 595 35723 14353 35728
rect 595 35689 624 35723
rect 658 35697 14289 35723
rect 658 35689 799 35697
rect 595 35663 799 35689
rect 833 35690 14289 35697
rect 833 35663 14114 35690
rect 595 35656 14114 35663
rect 14148 35689 14289 35690
rect 14323 35689 14353 35723
rect 14148 35656 14353 35689
rect 595 35655 14353 35656
rect 595 35621 624 35655
rect 658 35625 14289 35655
rect 658 35621 799 35625
rect 595 35591 799 35621
rect 833 35621 14289 35625
rect 14323 35621 14353 35655
rect 833 35618 14353 35621
rect 833 35591 14114 35618
rect 595 35587 14114 35591
rect 595 35553 624 35587
rect 658 35584 14114 35587
rect 14148 35587 14353 35618
rect 14148 35584 14289 35587
rect 658 35553 14289 35584
rect 14323 35553 14353 35587
rect 595 35519 799 35553
rect 833 35546 14353 35553
rect 833 35519 14114 35546
rect 595 35485 624 35519
rect 658 35512 14114 35519
rect 14148 35519 14353 35546
rect 14148 35512 14289 35519
rect 658 35485 14289 35512
rect 14323 35485 14353 35519
rect 595 35481 14353 35485
rect 595 35451 799 35481
rect 595 35417 624 35451
rect 658 35447 799 35451
rect 833 35474 14353 35481
rect 833 35447 14114 35474
rect 658 35440 14114 35447
rect 14148 35451 14353 35474
rect 14148 35440 14289 35451
rect 658 35417 14289 35440
rect 14323 35417 14353 35451
rect 595 35409 14353 35417
rect 595 35383 799 35409
rect 595 35349 624 35383
rect 658 35375 799 35383
rect 833 35402 14353 35409
rect 833 35375 14114 35402
rect 658 35368 14114 35375
rect 14148 35383 14353 35402
rect 14148 35368 14289 35383
rect 658 35349 14289 35368
rect 14323 35349 14353 35383
rect 595 35337 14353 35349
rect 595 35315 799 35337
rect 595 35281 624 35315
rect 658 35303 799 35315
rect 833 35330 14353 35337
rect 833 35303 14114 35330
rect 658 35296 14114 35303
rect 14148 35315 14353 35330
rect 14148 35296 14289 35315
rect 658 35281 14289 35296
rect 14323 35281 14353 35315
rect 595 35265 14353 35281
rect 595 35247 799 35265
rect 595 35213 624 35247
rect 658 35231 799 35247
rect 833 35258 14353 35265
rect 833 35231 14114 35258
rect 658 35224 14114 35231
rect 14148 35247 14353 35258
rect 14148 35224 14289 35247
rect 658 35213 14289 35224
rect 14323 35213 14353 35247
rect 595 35193 14353 35213
rect 595 35179 799 35193
rect 595 35145 624 35179
rect 658 35159 799 35179
rect 833 35186 14353 35193
rect 833 35159 14114 35186
rect 658 35152 14114 35159
rect 14148 35179 14353 35186
rect 14148 35152 14289 35179
rect 658 35145 14289 35152
rect 14323 35145 14353 35179
rect 595 35121 14353 35145
rect 595 35111 799 35121
rect 595 35077 624 35111
rect 658 35087 799 35111
rect 833 35114 14353 35121
rect 833 35087 14114 35114
rect 658 35080 14114 35087
rect 14148 35111 14353 35114
rect 14148 35080 14289 35111
rect 658 35077 14289 35080
rect 14323 35077 14353 35111
rect 595 35049 14353 35077
rect 595 35043 799 35049
rect 595 35009 624 35043
rect 658 35015 799 35043
rect 833 35043 14353 35049
rect 833 35042 14289 35043
rect 833 35015 14114 35042
rect 658 35009 14114 35015
rect 595 35008 14114 35009
rect 14148 35009 14289 35042
rect 14323 35009 14353 35043
rect 14148 35008 14353 35009
rect 595 34977 14353 35008
rect 595 34975 799 34977
rect 595 34941 624 34975
rect 658 34943 799 34975
rect 833 34975 14353 34977
rect 833 34970 14289 34975
rect 833 34943 14114 34970
rect 658 34941 14114 34943
rect 595 34936 14114 34941
rect 14148 34941 14289 34970
rect 14323 34941 14353 34975
rect 14148 34936 14353 34941
rect 595 34907 14353 34936
rect 595 34873 624 34907
rect 658 34905 14289 34907
rect 658 34873 799 34905
rect 595 34871 799 34873
rect 833 34898 14289 34905
rect 833 34871 14114 34898
rect 595 34864 14114 34871
rect 14148 34873 14289 34898
rect 14323 34873 14353 34907
rect 14148 34864 14353 34873
rect 595 34844 14353 34864
rect 595 34839 1018 34844
rect 595 34805 624 34839
rect 658 34833 1018 34839
rect 658 34805 799 34833
rect 595 34799 799 34805
rect 833 34799 1018 34833
rect 595 34771 1018 34799
rect 595 34737 624 34771
rect 658 34761 1018 34771
rect 658 34737 799 34761
rect 595 34727 799 34737
rect 833 34727 1018 34761
rect 13960 34839 14353 34844
rect 13960 34826 14289 34839
rect 13960 34792 14114 34826
rect 14148 34805 14289 34826
rect 14323 34805 14353 34839
rect 14148 34792 14353 34805
rect 13960 34771 14353 34792
rect 13960 34754 14289 34771
rect 595 34703 1018 34727
rect 595 34669 624 34703
rect 658 34689 1018 34703
rect 658 34669 799 34689
rect 595 34655 799 34669
rect 833 34655 1018 34689
rect 595 34635 1018 34655
rect 595 34601 624 34635
rect 658 34617 1018 34635
rect 658 34601 799 34617
rect 595 34583 799 34601
rect 833 34583 1018 34617
rect 595 34567 1018 34583
rect 595 34533 624 34567
rect 658 34545 1018 34567
rect 658 34533 799 34545
rect 595 34511 799 34533
rect 833 34511 1018 34545
rect 595 34499 1018 34511
rect 595 34465 624 34499
rect 658 34473 1018 34499
rect 658 34465 799 34473
rect 595 34439 799 34465
rect 833 34439 1018 34473
rect 595 34431 1018 34439
rect 595 34397 624 34431
rect 658 34401 1018 34431
rect 658 34397 799 34401
rect 595 34367 799 34397
rect 833 34367 1018 34401
rect 595 34363 1018 34367
rect 595 34329 624 34363
rect 658 34329 1018 34363
rect 595 34295 799 34329
rect 833 34295 1018 34329
rect 595 34261 624 34295
rect 658 34261 1018 34295
rect 595 34257 1018 34261
rect 595 34227 799 34257
rect 595 34193 624 34227
rect 658 34223 799 34227
rect 833 34223 1018 34257
rect 658 34193 1018 34223
rect 595 34185 1018 34193
rect 595 34159 799 34185
rect 595 34125 624 34159
rect 658 34151 799 34159
rect 833 34151 1018 34185
rect 658 34125 1018 34151
rect 595 34113 1018 34125
rect 595 34091 799 34113
rect 595 34057 624 34091
rect 658 34079 799 34091
rect 833 34079 1018 34113
rect 658 34057 1018 34079
rect 595 34041 1018 34057
rect 595 34023 799 34041
rect 595 33989 624 34023
rect 658 34007 799 34023
rect 833 34007 1018 34041
rect 658 33989 1018 34007
rect 595 33969 1018 33989
rect 595 33955 799 33969
rect 595 33921 624 33955
rect 658 33935 799 33955
rect 833 33935 1018 33969
rect 658 33921 1018 33935
rect 595 33897 1018 33921
rect 595 33887 799 33897
rect 595 33853 624 33887
rect 658 33863 799 33887
rect 833 33863 1018 33897
rect 658 33853 1018 33863
rect 595 33825 1018 33853
rect 595 33819 799 33825
rect 595 33785 624 33819
rect 658 33791 799 33819
rect 833 33791 1018 33825
rect 658 33785 1018 33791
rect 595 33753 1018 33785
rect 595 33751 799 33753
rect 595 33717 624 33751
rect 658 33719 799 33751
rect 833 33719 1018 33753
rect 658 33717 1018 33719
rect 595 33683 1018 33717
rect 595 33649 624 33683
rect 658 33681 1018 33683
rect 658 33649 799 33681
rect 595 33647 799 33649
rect 833 33647 1018 33681
rect 595 33615 1018 33647
rect 595 33581 624 33615
rect 658 33609 1018 33615
rect 658 33581 799 33609
rect 595 33575 799 33581
rect 833 33575 1018 33609
rect 595 33547 1018 33575
rect 595 33513 624 33547
rect 658 33537 1018 33547
rect 658 33513 799 33537
rect 595 33503 799 33513
rect 833 33503 1018 33537
rect 595 33479 1018 33503
rect 595 33445 624 33479
rect 658 33465 1018 33479
rect 658 33445 799 33465
rect 595 33431 799 33445
rect 833 33431 1018 33465
rect 595 33411 1018 33431
rect 595 33377 624 33411
rect 658 33393 1018 33411
rect 658 33377 799 33393
rect 595 33359 799 33377
rect 833 33359 1018 33393
rect 595 33343 1018 33359
rect 595 33309 624 33343
rect 658 33321 1018 33343
rect 658 33309 799 33321
rect 595 33287 799 33309
rect 833 33287 1018 33321
rect 595 33275 1018 33287
rect 595 33241 624 33275
rect 658 33249 1018 33275
rect 658 33241 799 33249
rect 595 33215 799 33241
rect 833 33215 1018 33249
rect 595 33207 1018 33215
rect 595 33173 624 33207
rect 658 33177 1018 33207
rect 658 33173 799 33177
rect 595 33143 799 33173
rect 833 33143 1018 33177
rect 595 33139 1018 33143
rect 595 33105 624 33139
rect 658 33105 1018 33139
rect 595 33071 799 33105
rect 833 33071 1018 33105
rect 595 33037 624 33071
rect 658 33037 1018 33071
rect 595 33033 1018 33037
rect 595 33003 799 33033
rect 595 32969 624 33003
rect 658 32999 799 33003
rect 833 32999 1018 33033
rect 658 32969 1018 32999
rect 595 32961 1018 32969
rect 595 32935 799 32961
rect 595 32901 624 32935
rect 658 32927 799 32935
rect 833 32927 1018 32961
rect 658 32901 1018 32927
rect 595 32889 1018 32901
rect 595 32867 799 32889
rect 595 32833 624 32867
rect 658 32855 799 32867
rect 833 32855 1018 32889
rect 658 32833 1018 32855
rect 595 32817 1018 32833
rect 595 32799 799 32817
rect 595 32765 624 32799
rect 658 32783 799 32799
rect 833 32783 1018 32817
rect 658 32765 1018 32783
rect 595 32745 1018 32765
rect 595 32731 799 32745
rect 595 32697 624 32731
rect 658 32711 799 32731
rect 833 32711 1018 32745
rect 658 32697 1018 32711
rect 595 32673 1018 32697
rect 595 32663 799 32673
rect 595 32629 624 32663
rect 658 32639 799 32663
rect 833 32639 1018 32673
rect 658 32629 1018 32639
rect 595 32601 1018 32629
rect 595 32595 799 32601
rect 595 32561 624 32595
rect 658 32567 799 32595
rect 833 32567 1018 32601
rect 658 32561 1018 32567
rect 595 32529 1018 32561
rect 595 32527 799 32529
rect 595 32493 624 32527
rect 658 32495 799 32527
rect 833 32495 1018 32529
rect 658 32493 1018 32495
rect 595 32459 1018 32493
rect 595 32425 624 32459
rect 658 32457 1018 32459
rect 658 32425 799 32457
rect 595 32423 799 32425
rect 833 32423 1018 32457
rect 595 32391 1018 32423
rect 595 32357 624 32391
rect 658 32385 1018 32391
rect 658 32357 799 32385
rect 595 32351 799 32357
rect 833 32351 1018 32385
rect 595 32323 1018 32351
rect 595 32289 624 32323
rect 658 32313 1018 32323
rect 658 32289 799 32313
rect 595 32279 799 32289
rect 833 32279 1018 32313
rect 595 32255 1018 32279
rect 595 32221 624 32255
rect 658 32241 1018 32255
rect 658 32221 799 32241
rect 595 32207 799 32221
rect 833 32207 1018 32241
rect 595 32187 1018 32207
rect 595 32153 624 32187
rect 658 32169 1018 32187
rect 658 32153 799 32169
rect 595 32135 799 32153
rect 833 32135 1018 32169
rect 595 32119 1018 32135
rect 595 32085 624 32119
rect 658 32097 1018 32119
rect 658 32085 799 32097
rect 595 32063 799 32085
rect 833 32063 1018 32097
rect 595 32051 1018 32063
rect 595 32017 624 32051
rect 658 32025 1018 32051
rect 658 32017 799 32025
rect 595 31991 799 32017
rect 833 31991 1018 32025
rect 595 31983 1018 31991
rect 595 31949 624 31983
rect 658 31953 1018 31983
rect 658 31949 799 31953
rect 595 31919 799 31949
rect 833 31919 1018 31953
rect 595 31915 1018 31919
rect 595 31881 624 31915
rect 658 31881 1018 31915
rect 595 31847 799 31881
rect 833 31847 1018 31881
rect 595 31813 624 31847
rect 658 31813 1018 31847
rect 595 31809 1018 31813
rect 595 31779 799 31809
rect 595 31745 624 31779
rect 658 31775 799 31779
rect 833 31775 1018 31809
rect 658 31745 1018 31775
rect 595 31737 1018 31745
rect 595 31711 799 31737
rect 595 31677 624 31711
rect 658 31703 799 31711
rect 833 31703 1018 31737
rect 658 31677 1018 31703
rect 595 31665 1018 31677
rect 595 31643 799 31665
rect 595 31609 624 31643
rect 658 31631 799 31643
rect 833 31631 1018 31665
rect 658 31609 1018 31631
rect 595 31593 1018 31609
rect 595 31575 799 31593
rect 595 31541 624 31575
rect 658 31559 799 31575
rect 833 31559 1018 31593
rect 658 31541 1018 31559
rect 595 31521 1018 31541
rect 595 31507 799 31521
rect 595 31473 624 31507
rect 658 31487 799 31507
rect 833 31487 1018 31521
rect 658 31473 1018 31487
rect 595 31449 1018 31473
rect 595 31439 799 31449
rect 595 31405 624 31439
rect 658 31415 799 31439
rect 833 31415 1018 31449
rect 658 31405 1018 31415
rect 595 31377 1018 31405
rect 595 31371 799 31377
rect 595 31337 624 31371
rect 658 31343 799 31371
rect 833 31343 1018 31377
rect 658 31337 1018 31343
rect 595 31305 1018 31337
rect 595 31303 799 31305
rect 595 31269 624 31303
rect 658 31271 799 31303
rect 833 31271 1018 31305
rect 658 31269 1018 31271
rect 595 31235 1018 31269
rect 595 31201 624 31235
rect 658 31233 1018 31235
rect 658 31201 799 31233
rect 595 31199 799 31201
rect 833 31199 1018 31233
rect 595 31167 1018 31199
rect 595 31133 624 31167
rect 658 31161 1018 31167
rect 658 31133 799 31161
rect 595 31127 799 31133
rect 833 31127 1018 31161
rect 595 31099 1018 31127
rect 595 31065 624 31099
rect 658 31089 1018 31099
rect 658 31065 799 31089
rect 595 31055 799 31065
rect 833 31055 1018 31089
rect 595 31031 1018 31055
rect 595 30997 624 31031
rect 658 31017 1018 31031
rect 658 30997 799 31017
rect 595 30983 799 30997
rect 833 30983 1018 31017
rect 595 30963 1018 30983
rect 595 30929 624 30963
rect 658 30945 1018 30963
rect 658 30929 799 30945
rect 595 30911 799 30929
rect 833 30911 1018 30945
rect 595 30895 1018 30911
rect 595 30861 624 30895
rect 658 30873 1018 30895
rect 658 30861 799 30873
rect 595 30839 799 30861
rect 833 30839 1018 30873
rect 595 30827 1018 30839
rect 595 30793 624 30827
rect 658 30801 1018 30827
rect 658 30793 799 30801
rect 595 30767 799 30793
rect 833 30767 1018 30801
rect 595 30759 1018 30767
rect 595 30725 624 30759
rect 658 30729 1018 30759
rect 658 30725 799 30729
rect 595 30695 799 30725
rect 833 30695 1018 30729
rect 595 30691 1018 30695
rect 595 30657 624 30691
rect 658 30657 1018 30691
rect 595 30623 799 30657
rect 833 30623 1018 30657
rect 595 30589 624 30623
rect 658 30589 1018 30623
rect 595 30585 1018 30589
rect 595 30555 799 30585
rect 595 30521 624 30555
rect 658 30551 799 30555
rect 833 30551 1018 30585
rect 658 30521 1018 30551
rect 595 30513 1018 30521
rect 595 30487 799 30513
rect 595 30453 624 30487
rect 658 30479 799 30487
rect 833 30479 1018 30513
rect 658 30453 1018 30479
rect 595 30441 1018 30453
rect 595 30419 799 30441
rect 595 30385 624 30419
rect 658 30407 799 30419
rect 833 30407 1018 30441
rect 658 30385 1018 30407
rect 595 30369 1018 30385
rect 595 30351 799 30369
rect 595 30317 624 30351
rect 658 30335 799 30351
rect 833 30335 1018 30369
rect 658 30317 1018 30335
rect 595 30297 1018 30317
rect 595 30283 799 30297
rect 595 30249 624 30283
rect 658 30263 799 30283
rect 833 30263 1018 30297
rect 658 30249 1018 30263
rect 595 30225 1018 30249
rect 595 30215 799 30225
rect 595 30181 624 30215
rect 658 30191 799 30215
rect 833 30191 1018 30225
rect 658 30181 1018 30191
rect 595 30153 1018 30181
rect 595 30147 799 30153
rect 595 30113 624 30147
rect 658 30119 799 30147
rect 833 30119 1018 30153
rect 658 30113 1018 30119
rect 595 30081 1018 30113
rect 595 30079 799 30081
rect 595 30045 624 30079
rect 658 30047 799 30079
rect 833 30047 1018 30081
rect 658 30045 1018 30047
rect 595 30011 1018 30045
rect 595 29977 624 30011
rect 658 30009 1018 30011
rect 658 29977 799 30009
rect 595 29975 799 29977
rect 833 29975 1018 30009
rect 595 29943 1018 29975
rect 595 29909 624 29943
rect 658 29937 1018 29943
rect 658 29909 799 29937
rect 595 29903 799 29909
rect 833 29903 1018 29937
rect 595 29875 1018 29903
rect 595 29841 624 29875
rect 658 29865 1018 29875
rect 658 29841 799 29865
rect 595 29831 799 29841
rect 833 29831 1018 29865
rect 595 29807 1018 29831
rect 595 29773 624 29807
rect 658 29793 1018 29807
rect 658 29773 799 29793
rect 595 29759 799 29773
rect 833 29759 1018 29793
rect 595 29739 1018 29759
rect 595 29705 624 29739
rect 658 29721 1018 29739
rect 658 29705 799 29721
rect 595 29687 799 29705
rect 833 29687 1018 29721
rect 595 29671 1018 29687
rect 595 29637 624 29671
rect 658 29649 1018 29671
rect 658 29637 799 29649
rect 595 29615 799 29637
rect 833 29615 1018 29649
rect 595 29603 1018 29615
rect 595 29569 624 29603
rect 658 29577 1018 29603
rect 658 29569 799 29577
rect 595 29543 799 29569
rect 833 29543 1018 29577
rect 595 29535 1018 29543
rect 595 29501 624 29535
rect 658 29505 1018 29535
rect 658 29501 799 29505
rect 595 29471 799 29501
rect 833 29471 1018 29505
rect 595 29467 1018 29471
rect 595 29433 624 29467
rect 658 29433 1018 29467
rect 595 29399 799 29433
rect 833 29399 1018 29433
rect 595 29365 624 29399
rect 658 29365 1018 29399
rect 595 29361 1018 29365
rect 595 29331 799 29361
rect 595 29297 624 29331
rect 658 29327 799 29331
rect 833 29327 1018 29361
rect 658 29297 1018 29327
rect 595 29289 1018 29297
rect 595 29263 799 29289
rect 595 29229 624 29263
rect 658 29255 799 29263
rect 833 29255 1018 29289
rect 658 29229 1018 29255
rect 595 29217 1018 29229
rect 595 29195 799 29217
rect 595 29161 624 29195
rect 658 29183 799 29195
rect 833 29183 1018 29217
rect 658 29161 1018 29183
rect 595 29145 1018 29161
rect 595 29127 799 29145
rect 595 29093 624 29127
rect 658 29111 799 29127
rect 833 29111 1018 29145
rect 658 29093 1018 29111
rect 595 29073 1018 29093
rect 595 29059 799 29073
rect 595 29025 624 29059
rect 658 29039 799 29059
rect 833 29039 1018 29073
rect 658 29025 1018 29039
rect 595 29001 1018 29025
rect 595 28991 799 29001
rect 595 28957 624 28991
rect 658 28967 799 28991
rect 833 28967 1018 29001
rect 658 28957 1018 28967
rect 595 28929 1018 28957
rect 595 28923 799 28929
rect 595 28889 624 28923
rect 658 28895 799 28923
rect 833 28895 1018 28929
rect 658 28889 1018 28895
rect 595 28857 1018 28889
rect 595 28855 799 28857
rect 595 28821 624 28855
rect 658 28823 799 28855
rect 833 28823 1018 28857
rect 658 28821 1018 28823
rect 595 28787 1018 28821
rect 595 28753 624 28787
rect 658 28785 1018 28787
rect 658 28753 799 28785
rect 595 28751 799 28753
rect 833 28751 1018 28785
rect 595 28719 1018 28751
rect 595 28685 624 28719
rect 658 28713 1018 28719
rect 658 28685 799 28713
rect 595 28679 799 28685
rect 833 28679 1018 28713
rect 595 28651 1018 28679
rect 595 28617 624 28651
rect 658 28641 1018 28651
rect 658 28617 799 28641
rect 595 28607 799 28617
rect 833 28607 1018 28641
rect 595 28583 1018 28607
rect 595 28549 624 28583
rect 658 28569 1018 28583
rect 658 28549 799 28569
rect 595 28535 799 28549
rect 833 28535 1018 28569
rect 595 28515 1018 28535
rect 595 28481 624 28515
rect 658 28497 1018 28515
rect 658 28481 799 28497
rect 595 28463 799 28481
rect 833 28463 1018 28497
rect 595 28447 1018 28463
rect 595 28413 624 28447
rect 658 28425 1018 28447
rect 658 28413 799 28425
rect 595 28391 799 28413
rect 833 28391 1018 28425
rect 595 28379 1018 28391
rect 595 28345 624 28379
rect 658 28353 1018 28379
rect 658 28345 799 28353
rect 595 28319 799 28345
rect 833 28319 1018 28353
rect 595 28311 1018 28319
rect 595 28277 624 28311
rect 658 28281 1018 28311
rect 658 28277 799 28281
rect 595 28247 799 28277
rect 833 28247 1018 28281
rect 595 28243 1018 28247
rect 595 28209 624 28243
rect 658 28209 1018 28243
rect 595 28175 799 28209
rect 833 28175 1018 28209
rect 595 28141 624 28175
rect 658 28141 1018 28175
rect 595 28137 1018 28141
rect 595 28107 799 28137
rect 595 28073 624 28107
rect 658 28103 799 28107
rect 833 28103 1018 28137
rect 658 28073 1018 28103
rect 595 28065 1018 28073
rect 595 28039 799 28065
rect 595 28005 624 28039
rect 658 28031 799 28039
rect 833 28031 1018 28065
rect 658 28005 1018 28031
rect 595 27993 1018 28005
rect 595 27971 799 27993
rect 595 27937 624 27971
rect 658 27959 799 27971
rect 833 27959 1018 27993
rect 658 27937 1018 27959
rect 595 27921 1018 27937
rect 595 27903 799 27921
rect 595 27869 624 27903
rect 658 27887 799 27903
rect 833 27887 1018 27921
rect 658 27869 1018 27887
rect 595 27849 1018 27869
rect 595 27835 799 27849
rect 595 27801 624 27835
rect 658 27815 799 27835
rect 833 27815 1018 27849
rect 658 27801 1018 27815
rect 595 27777 1018 27801
rect 595 27767 799 27777
rect 595 27733 624 27767
rect 658 27743 799 27767
rect 833 27743 1018 27777
rect 658 27733 1018 27743
rect 595 27705 1018 27733
rect 595 27699 799 27705
rect 595 27665 624 27699
rect 658 27671 799 27699
rect 833 27671 1018 27705
rect 658 27665 1018 27671
rect 595 27633 1018 27665
rect 595 27631 799 27633
rect 595 27597 624 27631
rect 658 27599 799 27631
rect 833 27599 1018 27633
rect 658 27597 1018 27599
rect 595 27563 1018 27597
rect 595 27529 624 27563
rect 658 27561 1018 27563
rect 658 27529 799 27561
rect 595 27527 799 27529
rect 833 27527 1018 27561
rect 595 27495 1018 27527
rect 595 27461 624 27495
rect 658 27489 1018 27495
rect 658 27461 799 27489
rect 595 27455 799 27461
rect 833 27455 1018 27489
rect 595 27427 1018 27455
rect 595 27393 624 27427
rect 658 27417 1018 27427
rect 658 27393 799 27417
rect 595 27383 799 27393
rect 833 27383 1018 27417
rect 595 27359 1018 27383
rect 595 27325 624 27359
rect 658 27345 1018 27359
rect 658 27325 799 27345
rect 595 27311 799 27325
rect 833 27311 1018 27345
rect 595 27291 1018 27311
rect 595 27257 624 27291
rect 658 27273 1018 27291
rect 658 27257 799 27273
rect 595 27239 799 27257
rect 833 27239 1018 27273
rect 595 27223 1018 27239
rect 595 27189 624 27223
rect 658 27201 1018 27223
rect 658 27189 799 27201
rect 595 27167 799 27189
rect 833 27167 1018 27201
rect 595 27155 1018 27167
rect 595 27121 624 27155
rect 658 27129 1018 27155
rect 658 27121 799 27129
rect 595 27095 799 27121
rect 833 27095 1018 27129
rect 595 27087 1018 27095
rect 595 27053 624 27087
rect 658 27057 1018 27087
rect 658 27053 799 27057
rect 595 27023 799 27053
rect 833 27023 1018 27057
rect 595 27019 1018 27023
rect 595 26985 624 27019
rect 658 26985 1018 27019
rect 595 26951 799 26985
rect 833 26951 1018 26985
rect 595 26917 624 26951
rect 658 26917 1018 26951
rect 595 26913 1018 26917
rect 595 26883 799 26913
rect 595 26849 624 26883
rect 658 26879 799 26883
rect 833 26879 1018 26913
rect 658 26849 1018 26879
rect 595 26841 1018 26849
rect 595 26815 799 26841
rect 595 26781 624 26815
rect 658 26807 799 26815
rect 833 26807 1018 26841
rect 658 26781 1018 26807
rect 595 26769 1018 26781
rect 595 26747 799 26769
rect 595 26713 624 26747
rect 658 26735 799 26747
rect 833 26735 1018 26769
rect 658 26713 1018 26735
rect 595 26697 1018 26713
rect 595 26679 799 26697
rect 595 26645 624 26679
rect 658 26663 799 26679
rect 833 26663 1018 26697
rect 658 26645 1018 26663
rect 595 26625 1018 26645
rect 595 26611 799 26625
rect 595 26577 624 26611
rect 658 26591 799 26611
rect 833 26591 1018 26625
rect 658 26577 1018 26591
rect 595 26553 1018 26577
rect 595 26543 799 26553
rect 595 26509 624 26543
rect 658 26519 799 26543
rect 833 26519 1018 26553
rect 658 26509 1018 26519
rect 595 26481 1018 26509
rect 595 26475 799 26481
rect 595 26441 624 26475
rect 658 26447 799 26475
rect 833 26447 1018 26481
rect 658 26441 1018 26447
rect 595 26409 1018 26441
rect 595 26407 799 26409
rect 595 26373 624 26407
rect 658 26375 799 26407
rect 833 26375 1018 26409
rect 658 26373 1018 26375
rect 595 26339 1018 26373
rect 595 26305 624 26339
rect 658 26337 1018 26339
rect 658 26305 799 26337
rect 595 26303 799 26305
rect 833 26303 1018 26337
rect 595 26271 1018 26303
rect 595 26237 624 26271
rect 658 26265 1018 26271
rect 658 26237 799 26265
rect 595 26231 799 26237
rect 833 26231 1018 26265
rect 595 26203 1018 26231
rect 595 26169 624 26203
rect 658 26193 1018 26203
rect 658 26169 799 26193
rect 595 26159 799 26169
rect 833 26159 1018 26193
rect 595 26135 1018 26159
rect 595 26101 624 26135
rect 658 26121 1018 26135
rect 658 26101 799 26121
rect 595 26087 799 26101
rect 833 26087 1018 26121
rect 595 26067 1018 26087
rect 595 26033 624 26067
rect 658 26049 1018 26067
rect 658 26033 799 26049
rect 595 26015 799 26033
rect 833 26015 1018 26049
rect 595 25999 1018 26015
rect 595 25965 624 25999
rect 658 25977 1018 25999
rect 658 25965 799 25977
rect 595 25943 799 25965
rect 833 25943 1018 25977
rect 595 25931 1018 25943
rect 595 25897 624 25931
rect 658 25905 1018 25931
rect 658 25897 799 25905
rect 595 25871 799 25897
rect 833 25871 1018 25905
rect 595 25863 1018 25871
rect 595 25829 624 25863
rect 658 25833 1018 25863
rect 658 25829 799 25833
rect 595 25799 799 25829
rect 833 25799 1018 25833
rect 595 25795 1018 25799
rect 595 25761 624 25795
rect 658 25761 1018 25795
rect 595 25727 799 25761
rect 833 25727 1018 25761
rect 595 25693 624 25727
rect 658 25693 1018 25727
rect 595 25689 1018 25693
rect 595 25659 799 25689
rect 595 25625 624 25659
rect 658 25655 799 25659
rect 833 25655 1018 25689
rect 658 25625 1018 25655
rect 595 25617 1018 25625
rect 595 25591 799 25617
rect 595 25557 624 25591
rect 658 25583 799 25591
rect 833 25583 1018 25617
rect 658 25557 1018 25583
rect 595 25545 1018 25557
rect 595 25523 799 25545
rect 595 25489 624 25523
rect 658 25511 799 25523
rect 833 25511 1018 25545
rect 658 25489 1018 25511
rect 595 25473 1018 25489
rect 595 25455 799 25473
rect 595 25421 624 25455
rect 658 25439 799 25455
rect 833 25439 1018 25473
rect 658 25421 1018 25439
rect 595 25401 1018 25421
rect 595 25387 799 25401
rect 595 25353 624 25387
rect 658 25367 799 25387
rect 833 25367 1018 25401
rect 658 25353 1018 25367
rect 595 25329 1018 25353
rect 595 25319 799 25329
rect 595 25285 624 25319
rect 658 25295 799 25319
rect 833 25295 1018 25329
rect 658 25285 1018 25295
rect 595 25257 1018 25285
rect 595 25251 799 25257
rect 595 25217 624 25251
rect 658 25223 799 25251
rect 833 25223 1018 25257
rect 658 25217 1018 25223
rect 595 25185 1018 25217
rect 595 25183 799 25185
rect 595 25149 624 25183
rect 658 25151 799 25183
rect 833 25151 1018 25185
rect 658 25149 1018 25151
rect 595 25115 1018 25149
rect 595 25081 624 25115
rect 658 25113 1018 25115
rect 658 25081 799 25113
rect 595 25079 799 25081
rect 833 25079 1018 25113
rect 595 25047 1018 25079
rect 595 25013 624 25047
rect 658 25041 1018 25047
rect 658 25013 799 25041
rect 595 25007 799 25013
rect 833 25007 1018 25041
rect 595 24979 1018 25007
rect 595 24945 624 24979
rect 658 24969 1018 24979
rect 658 24945 799 24969
rect 595 24935 799 24945
rect 833 24935 1018 24969
rect 595 24911 1018 24935
rect 595 24877 624 24911
rect 658 24897 1018 24911
rect 658 24877 799 24897
rect 595 24863 799 24877
rect 833 24863 1018 24897
rect 595 24843 1018 24863
rect 595 24809 624 24843
rect 658 24825 1018 24843
rect 658 24809 799 24825
rect 595 24791 799 24809
rect 833 24791 1018 24825
rect 595 24775 1018 24791
rect 595 24741 624 24775
rect 658 24753 1018 24775
rect 658 24741 799 24753
rect 595 24719 799 24741
rect 833 24719 1018 24753
rect 595 24707 1018 24719
rect 595 24673 624 24707
rect 658 24681 1018 24707
rect 658 24673 799 24681
rect 595 24647 799 24673
rect 833 24647 1018 24681
rect 595 24639 1018 24647
rect 595 24605 624 24639
rect 658 24609 1018 24639
rect 658 24605 799 24609
rect 595 24575 799 24605
rect 833 24575 1018 24609
rect 595 24571 1018 24575
rect 595 24537 624 24571
rect 658 24537 1018 24571
rect 595 24503 799 24537
rect 833 24503 1018 24537
rect 595 24469 624 24503
rect 658 24469 1018 24503
rect 595 24465 1018 24469
rect 595 24435 799 24465
rect 595 24401 624 24435
rect 658 24431 799 24435
rect 833 24431 1018 24465
rect 658 24401 1018 24431
rect 595 24393 1018 24401
rect 595 24367 799 24393
rect 595 24333 624 24367
rect 658 24359 799 24367
rect 833 24359 1018 24393
rect 658 24333 1018 24359
rect 595 24321 1018 24333
rect 595 24299 799 24321
rect 595 24265 624 24299
rect 658 24287 799 24299
rect 833 24287 1018 24321
rect 658 24265 1018 24287
rect 595 24249 1018 24265
rect 595 24231 799 24249
rect 595 24197 624 24231
rect 658 24215 799 24231
rect 833 24215 1018 24249
rect 658 24197 1018 24215
rect 595 24177 1018 24197
rect 595 24163 799 24177
rect 595 24129 624 24163
rect 658 24143 799 24163
rect 833 24143 1018 24177
rect 658 24129 1018 24143
rect 595 24105 1018 24129
rect 595 24095 799 24105
rect 595 24061 624 24095
rect 658 24071 799 24095
rect 833 24071 1018 24105
rect 658 24061 1018 24071
rect 595 24033 1018 24061
rect 595 24027 799 24033
rect 595 23993 624 24027
rect 658 23999 799 24027
rect 833 23999 1018 24033
rect 658 23993 1018 23999
rect 595 23961 1018 23993
rect 595 23959 799 23961
rect 595 23925 624 23959
rect 658 23927 799 23959
rect 833 23927 1018 23961
rect 658 23925 1018 23927
rect 595 23891 1018 23925
rect 595 23857 624 23891
rect 658 23889 1018 23891
rect 658 23857 799 23889
rect 595 23855 799 23857
rect 833 23855 1018 23889
rect 595 23823 1018 23855
rect 595 23789 624 23823
rect 658 23817 1018 23823
rect 658 23789 799 23817
rect 595 23783 799 23789
rect 833 23783 1018 23817
rect 595 23755 1018 23783
rect 595 23721 624 23755
rect 658 23745 1018 23755
rect 658 23721 799 23745
rect 595 23711 799 23721
rect 833 23711 1018 23745
rect 595 23687 1018 23711
rect 595 23653 624 23687
rect 658 23673 1018 23687
rect 658 23653 799 23673
rect 595 23639 799 23653
rect 833 23639 1018 23673
rect 595 23619 1018 23639
rect 595 23585 624 23619
rect 658 23601 1018 23619
rect 658 23585 799 23601
rect 595 23567 799 23585
rect 833 23567 1018 23601
rect 595 23551 1018 23567
rect 595 23517 624 23551
rect 658 23529 1018 23551
rect 658 23517 799 23529
rect 595 23495 799 23517
rect 833 23495 1018 23529
rect 595 23483 1018 23495
rect 595 23449 624 23483
rect 658 23457 1018 23483
rect 658 23449 799 23457
rect 595 23423 799 23449
rect 833 23423 1018 23457
rect 595 23415 1018 23423
rect 595 23381 624 23415
rect 658 23385 1018 23415
rect 658 23381 799 23385
rect 595 23351 799 23381
rect 833 23351 1018 23385
rect 595 23347 1018 23351
rect 595 23313 624 23347
rect 658 23313 1018 23347
rect 595 23279 799 23313
rect 833 23279 1018 23313
rect 595 23245 624 23279
rect 658 23245 1018 23279
rect 595 23241 1018 23245
rect 595 23211 799 23241
rect 595 23177 624 23211
rect 658 23207 799 23211
rect 833 23207 1018 23241
rect 658 23177 1018 23207
rect 595 23169 1018 23177
rect 595 23143 799 23169
rect 595 23109 624 23143
rect 658 23135 799 23143
rect 833 23135 1018 23169
rect 658 23109 1018 23135
rect 595 23097 1018 23109
rect 595 23075 799 23097
rect 595 23041 624 23075
rect 658 23063 799 23075
rect 833 23063 1018 23097
rect 658 23041 1018 23063
rect 595 23025 1018 23041
rect 595 23007 799 23025
rect 595 22973 624 23007
rect 658 22991 799 23007
rect 833 22991 1018 23025
rect 658 22973 1018 22991
rect 595 22953 1018 22973
rect 595 22939 799 22953
rect 595 22905 624 22939
rect 658 22919 799 22939
rect 833 22919 1018 22953
rect 658 22905 1018 22919
rect 595 22881 1018 22905
rect 595 22871 799 22881
rect 595 22837 624 22871
rect 658 22847 799 22871
rect 833 22847 1018 22881
rect 658 22837 1018 22847
rect 595 22809 1018 22837
rect 595 22803 799 22809
rect 595 22769 624 22803
rect 658 22775 799 22803
rect 833 22775 1018 22809
rect 658 22769 1018 22775
rect 595 22737 1018 22769
rect 595 22735 799 22737
rect 595 22701 624 22735
rect 658 22703 799 22735
rect 833 22703 1018 22737
rect 658 22701 1018 22703
rect 595 22667 1018 22701
rect 595 22633 624 22667
rect 658 22665 1018 22667
rect 658 22633 799 22665
rect 595 22631 799 22633
rect 833 22631 1018 22665
rect 595 22599 1018 22631
rect 595 22565 624 22599
rect 658 22593 1018 22599
rect 658 22565 799 22593
rect 595 22559 799 22565
rect 833 22559 1018 22593
rect 595 22531 1018 22559
rect 595 22497 624 22531
rect 658 22521 1018 22531
rect 658 22497 799 22521
rect 595 22487 799 22497
rect 833 22487 1018 22521
rect 595 22463 1018 22487
rect 595 22429 624 22463
rect 658 22449 1018 22463
rect 658 22429 799 22449
rect 595 22415 799 22429
rect 833 22415 1018 22449
rect 595 22395 1018 22415
rect 595 22361 624 22395
rect 658 22377 1018 22395
rect 658 22361 799 22377
rect 595 22343 799 22361
rect 833 22343 1018 22377
rect 595 22327 1018 22343
rect 595 22293 624 22327
rect 658 22305 1018 22327
rect 658 22293 799 22305
rect 595 22271 799 22293
rect 833 22271 1018 22305
rect 595 22259 1018 22271
rect 595 22225 624 22259
rect 658 22233 1018 22259
rect 658 22225 799 22233
rect 595 22199 799 22225
rect 833 22199 1018 22233
rect 595 22191 1018 22199
rect 595 22157 624 22191
rect 658 22161 1018 22191
rect 658 22157 799 22161
rect 595 22127 799 22157
rect 833 22127 1018 22161
rect 595 22123 1018 22127
rect 595 22089 624 22123
rect 658 22089 1018 22123
rect 595 22055 799 22089
rect 833 22055 1018 22089
rect 595 22021 624 22055
rect 658 22021 1018 22055
rect 595 22017 1018 22021
rect 595 21987 799 22017
rect 595 21953 624 21987
rect 658 21983 799 21987
rect 833 21983 1018 22017
rect 658 21953 1018 21983
rect 595 21945 1018 21953
rect 595 21919 799 21945
rect 595 21885 624 21919
rect 658 21911 799 21919
rect 833 21911 1018 21945
rect 658 21885 1018 21911
rect 595 21873 1018 21885
rect 595 21851 799 21873
rect 595 21817 624 21851
rect 658 21839 799 21851
rect 833 21839 1018 21873
rect 658 21817 1018 21839
rect 595 21801 1018 21817
rect 595 21783 799 21801
rect 595 21749 624 21783
rect 658 21767 799 21783
rect 833 21767 1018 21801
rect 658 21749 1018 21767
rect 595 21729 1018 21749
rect 595 21715 799 21729
rect 595 21681 624 21715
rect 658 21695 799 21715
rect 833 21695 1018 21729
rect 658 21681 1018 21695
rect 595 21657 1018 21681
rect 595 21647 799 21657
rect 595 21613 624 21647
rect 658 21623 799 21647
rect 833 21623 1018 21657
rect 658 21613 1018 21623
rect 595 21585 1018 21613
rect 595 21579 799 21585
rect 595 21545 624 21579
rect 658 21551 799 21579
rect 833 21551 1018 21585
rect 658 21545 1018 21551
rect 595 21513 1018 21545
rect 595 21511 799 21513
rect 595 21477 624 21511
rect 658 21479 799 21511
rect 833 21479 1018 21513
rect 658 21477 1018 21479
rect 595 21443 1018 21477
rect 595 21409 624 21443
rect 658 21441 1018 21443
rect 658 21409 799 21441
rect 595 21407 799 21409
rect 833 21407 1018 21441
rect 595 21375 1018 21407
rect 595 21341 624 21375
rect 658 21369 1018 21375
rect 658 21341 799 21369
rect 595 21335 799 21341
rect 833 21335 1018 21369
rect 595 21307 1018 21335
rect 595 21273 624 21307
rect 658 21297 1018 21307
rect 658 21273 799 21297
rect 595 21263 799 21273
rect 833 21263 1018 21297
rect 595 21239 1018 21263
rect 595 21205 624 21239
rect 658 21225 1018 21239
rect 658 21205 799 21225
rect 595 21191 799 21205
rect 833 21191 1018 21225
rect 595 21171 1018 21191
rect 595 21137 624 21171
rect 658 21153 1018 21171
rect 658 21137 799 21153
rect 595 21119 799 21137
rect 833 21119 1018 21153
rect 595 21103 1018 21119
rect 595 21069 624 21103
rect 658 21081 1018 21103
rect 658 21069 799 21081
rect 595 21047 799 21069
rect 833 21047 1018 21081
rect 595 21035 1018 21047
rect 595 21001 624 21035
rect 658 21009 1018 21035
rect 658 21001 799 21009
rect 595 20975 799 21001
rect 833 20975 1018 21009
rect 595 20967 1018 20975
rect 595 20933 624 20967
rect 658 20937 1018 20967
rect 658 20933 799 20937
rect 595 20903 799 20933
rect 833 20903 1018 20937
rect 595 20899 1018 20903
rect 595 20865 624 20899
rect 658 20865 1018 20899
rect 595 20831 799 20865
rect 833 20831 1018 20865
rect 595 20797 624 20831
rect 658 20797 1018 20831
rect 595 20793 1018 20797
rect 595 20763 799 20793
rect 595 20729 624 20763
rect 658 20759 799 20763
rect 833 20759 1018 20793
rect 658 20729 1018 20759
rect 595 20721 1018 20729
rect 595 20695 799 20721
rect 595 20661 624 20695
rect 658 20687 799 20695
rect 833 20687 1018 20721
rect 658 20661 1018 20687
rect 595 20649 1018 20661
rect 595 20627 799 20649
rect 595 20593 624 20627
rect 658 20615 799 20627
rect 833 20615 1018 20649
rect 658 20593 1018 20615
rect 595 20577 1018 20593
rect 595 20559 799 20577
rect 595 20525 624 20559
rect 658 20543 799 20559
rect 833 20543 1018 20577
rect 658 20525 1018 20543
rect 595 20505 1018 20525
rect 595 20491 799 20505
rect 595 20457 624 20491
rect 658 20471 799 20491
rect 833 20471 1018 20505
rect 658 20457 1018 20471
rect 595 20433 1018 20457
rect 595 20423 799 20433
rect 595 20389 624 20423
rect 658 20399 799 20423
rect 833 20399 1018 20433
rect 658 20389 1018 20399
rect 595 20361 1018 20389
rect 595 20355 799 20361
rect 595 20321 624 20355
rect 658 20327 799 20355
rect 833 20327 1018 20361
rect 658 20321 1018 20327
rect 595 20289 1018 20321
rect 595 20287 799 20289
rect 595 20253 624 20287
rect 658 20255 799 20287
rect 833 20255 1018 20289
rect 658 20253 1018 20255
rect 595 20219 1018 20253
rect 595 20185 624 20219
rect 658 20217 1018 20219
rect 658 20185 799 20217
rect 595 20183 799 20185
rect 833 20183 1018 20217
rect 595 20151 1018 20183
rect 595 20117 624 20151
rect 658 20145 1018 20151
rect 658 20117 799 20145
rect 595 20111 799 20117
rect 833 20111 1018 20145
rect 595 20083 1018 20111
rect 595 20049 624 20083
rect 658 20073 1018 20083
rect 658 20049 799 20073
rect 595 20039 799 20049
rect 833 20039 1018 20073
rect 595 20015 1018 20039
rect 595 19981 624 20015
rect 658 20001 1018 20015
rect 658 19981 799 20001
rect 595 19967 799 19981
rect 833 19967 1018 20001
rect 595 19947 1018 19967
rect 595 19913 624 19947
rect 658 19929 1018 19947
rect 658 19913 799 19929
rect 595 19895 799 19913
rect 833 19895 1018 19929
rect 595 19879 1018 19895
rect 595 19845 624 19879
rect 658 19857 1018 19879
rect 658 19845 799 19857
rect 595 19823 799 19845
rect 833 19823 1018 19857
rect 595 19811 1018 19823
rect 595 19777 624 19811
rect 658 19785 1018 19811
rect 658 19777 799 19785
rect 595 19751 799 19777
rect 833 19751 1018 19785
rect 595 19743 1018 19751
rect 595 19709 624 19743
rect 658 19713 1018 19743
rect 658 19709 799 19713
rect 595 19679 799 19709
rect 833 19679 1018 19713
rect 595 19675 1018 19679
rect 595 19641 624 19675
rect 658 19641 1018 19675
rect 595 19607 799 19641
rect 833 19607 1018 19641
rect 595 19573 624 19607
rect 658 19573 1018 19607
rect 595 19569 1018 19573
rect 595 19539 799 19569
rect 595 19505 624 19539
rect 658 19535 799 19539
rect 833 19535 1018 19569
rect 658 19505 1018 19535
rect 595 19497 1018 19505
rect 595 19471 799 19497
rect 595 19437 624 19471
rect 658 19463 799 19471
rect 833 19463 1018 19497
rect 658 19437 1018 19463
rect 595 19425 1018 19437
rect 595 19403 799 19425
rect 595 19369 624 19403
rect 658 19391 799 19403
rect 833 19391 1018 19425
rect 658 19369 1018 19391
rect 595 19353 1018 19369
rect 595 19335 799 19353
rect 595 19301 624 19335
rect 658 19319 799 19335
rect 833 19319 1018 19353
rect 658 19301 1018 19319
rect 595 19281 1018 19301
rect 595 19267 799 19281
rect 595 19233 624 19267
rect 658 19247 799 19267
rect 833 19247 1018 19281
rect 658 19233 1018 19247
rect 595 19209 1018 19233
rect 595 19199 799 19209
rect 595 19165 624 19199
rect 658 19175 799 19199
rect 833 19175 1018 19209
rect 658 19165 1018 19175
rect 595 19137 1018 19165
rect 595 19131 799 19137
rect 595 19097 624 19131
rect 658 19103 799 19131
rect 833 19103 1018 19137
rect 658 19097 1018 19103
rect 595 19065 1018 19097
rect 595 19063 799 19065
rect 595 19029 624 19063
rect 658 19031 799 19063
rect 833 19031 1018 19065
rect 658 19029 1018 19031
rect 595 18995 1018 19029
rect 595 18961 624 18995
rect 658 18993 1018 18995
rect 658 18961 799 18993
rect 595 18959 799 18961
rect 833 18959 1018 18993
rect 595 18927 1018 18959
rect 595 18893 624 18927
rect 658 18921 1018 18927
rect 658 18893 799 18921
rect 595 18887 799 18893
rect 833 18887 1018 18921
rect 595 18859 1018 18887
rect 595 18825 624 18859
rect 658 18849 1018 18859
rect 658 18825 799 18849
rect 595 18815 799 18825
rect 833 18815 1018 18849
rect 595 18791 1018 18815
rect 595 18757 624 18791
rect 658 18777 1018 18791
rect 658 18757 799 18777
rect 595 18743 799 18757
rect 833 18743 1018 18777
rect 595 18723 1018 18743
rect 595 18689 624 18723
rect 658 18705 1018 18723
rect 658 18689 799 18705
rect 595 18671 799 18689
rect 833 18671 1018 18705
rect 595 18655 1018 18671
rect 595 18621 624 18655
rect 658 18633 1018 18655
rect 658 18621 799 18633
rect 595 18599 799 18621
rect 833 18599 1018 18633
rect 595 18587 1018 18599
rect 595 18553 624 18587
rect 658 18561 1018 18587
rect 658 18553 799 18561
rect 595 18527 799 18553
rect 833 18527 1018 18561
rect 595 18519 1018 18527
rect 595 18485 624 18519
rect 658 18489 1018 18519
rect 658 18485 799 18489
rect 595 18455 799 18485
rect 833 18455 1018 18489
rect 595 18451 1018 18455
rect 595 18417 624 18451
rect 658 18417 1018 18451
rect 595 18383 799 18417
rect 833 18383 1018 18417
rect 595 18349 624 18383
rect 658 18349 1018 18383
rect 595 18345 1018 18349
rect 595 18315 799 18345
rect 595 18281 624 18315
rect 658 18311 799 18315
rect 833 18311 1018 18345
rect 658 18281 1018 18311
rect 595 18273 1018 18281
rect 595 18247 799 18273
rect 595 18213 624 18247
rect 658 18239 799 18247
rect 833 18239 1018 18273
rect 658 18213 1018 18239
rect 595 18201 1018 18213
rect 595 18179 799 18201
rect 595 18145 624 18179
rect 658 18167 799 18179
rect 833 18167 1018 18201
rect 658 18145 1018 18167
rect 595 18129 1018 18145
rect 595 18111 799 18129
rect 595 18077 624 18111
rect 658 18095 799 18111
rect 833 18095 1018 18129
rect 658 18077 1018 18095
rect 595 18057 1018 18077
rect 595 18043 799 18057
rect 595 18009 624 18043
rect 658 18023 799 18043
rect 833 18023 1018 18057
rect 658 18009 1018 18023
rect 595 17985 1018 18009
rect 595 17975 799 17985
rect 595 17941 624 17975
rect 658 17951 799 17975
rect 833 17951 1018 17985
rect 658 17941 1018 17951
rect 595 17913 1018 17941
rect 595 17907 799 17913
rect 595 17873 624 17907
rect 658 17879 799 17907
rect 833 17879 1018 17913
rect 658 17873 1018 17879
rect 595 17841 1018 17873
rect 595 17839 799 17841
rect 595 17805 624 17839
rect 658 17807 799 17839
rect 833 17807 1018 17841
rect 658 17805 1018 17807
rect 595 17771 1018 17805
rect 595 17737 624 17771
rect 658 17769 1018 17771
rect 658 17737 799 17769
rect 595 17735 799 17737
rect 833 17735 1018 17769
rect 595 17703 1018 17735
rect 595 17669 624 17703
rect 658 17697 1018 17703
rect 658 17669 799 17697
rect 595 17663 799 17669
rect 833 17663 1018 17697
rect 595 17635 1018 17663
rect 595 17601 624 17635
rect 658 17625 1018 17635
rect 658 17601 799 17625
rect 595 17591 799 17601
rect 833 17591 1018 17625
rect 595 17567 1018 17591
rect 595 17533 624 17567
rect 658 17553 1018 17567
rect 658 17533 799 17553
rect 595 17519 799 17533
rect 833 17519 1018 17553
rect 595 17499 1018 17519
rect 595 17465 624 17499
rect 658 17481 1018 17499
rect 658 17465 799 17481
rect 595 17447 799 17465
rect 833 17447 1018 17481
rect 595 17431 1018 17447
rect 595 17397 624 17431
rect 658 17409 1018 17431
rect 658 17397 799 17409
rect 595 17375 799 17397
rect 833 17375 1018 17409
rect 595 17363 1018 17375
rect 595 17329 624 17363
rect 658 17337 1018 17363
rect 658 17329 799 17337
rect 595 17303 799 17329
rect 833 17303 1018 17337
rect 595 17295 1018 17303
rect 595 17261 624 17295
rect 658 17265 1018 17295
rect 658 17261 799 17265
rect 595 17231 799 17261
rect 833 17231 1018 17265
rect 595 17227 1018 17231
rect 595 17193 624 17227
rect 658 17193 1018 17227
rect 595 17159 799 17193
rect 833 17159 1018 17193
rect 595 17125 624 17159
rect 658 17125 1018 17159
rect 595 17121 1018 17125
rect 595 17091 799 17121
rect 595 17057 624 17091
rect 658 17087 799 17091
rect 833 17087 1018 17121
rect 658 17057 1018 17087
rect 595 17049 1018 17057
rect 595 17023 799 17049
rect 595 16989 624 17023
rect 658 17015 799 17023
rect 833 17015 1018 17049
rect 658 16989 1018 17015
rect 595 16977 1018 16989
rect 595 16955 799 16977
rect 595 16921 624 16955
rect 658 16943 799 16955
rect 833 16943 1018 16977
rect 658 16921 1018 16943
rect 595 16905 1018 16921
rect 595 16887 799 16905
rect 595 16853 624 16887
rect 658 16871 799 16887
rect 833 16871 1018 16905
rect 658 16853 1018 16871
rect 595 16833 1018 16853
rect 595 16819 799 16833
rect 595 16785 624 16819
rect 658 16799 799 16819
rect 833 16799 1018 16833
rect 658 16785 1018 16799
rect 595 16761 1018 16785
rect 595 16751 799 16761
rect 595 16717 624 16751
rect 658 16727 799 16751
rect 833 16727 1018 16761
rect 658 16717 1018 16727
rect 595 16689 1018 16717
rect 595 16683 799 16689
rect 595 16649 624 16683
rect 658 16655 799 16683
rect 833 16655 1018 16689
rect 658 16649 1018 16655
rect 595 16617 1018 16649
rect 595 16615 799 16617
rect 595 16581 624 16615
rect 658 16583 799 16615
rect 833 16583 1018 16617
rect 658 16581 1018 16583
rect 595 16547 1018 16581
rect 595 16513 624 16547
rect 658 16545 1018 16547
rect 658 16513 799 16545
rect 595 16511 799 16513
rect 833 16511 1018 16545
rect 595 16479 1018 16511
rect 595 16445 624 16479
rect 658 16473 1018 16479
rect 658 16445 799 16473
rect 595 16439 799 16445
rect 833 16439 1018 16473
rect 595 16411 1018 16439
rect 595 16377 624 16411
rect 658 16401 1018 16411
rect 658 16377 799 16401
rect 595 16367 799 16377
rect 833 16367 1018 16401
rect 595 16343 1018 16367
rect 595 16309 624 16343
rect 658 16329 1018 16343
rect 658 16309 799 16329
rect 595 16295 799 16309
rect 833 16295 1018 16329
rect 595 16275 1018 16295
rect 595 16241 624 16275
rect 658 16257 1018 16275
rect 658 16241 799 16257
rect 595 16223 799 16241
rect 833 16223 1018 16257
rect 595 16207 1018 16223
rect 595 16173 624 16207
rect 658 16185 1018 16207
rect 658 16173 799 16185
rect 595 16151 799 16173
rect 833 16151 1018 16185
rect 595 16139 1018 16151
rect 595 16105 624 16139
rect 658 16113 1018 16139
rect 658 16105 799 16113
rect 595 16079 799 16105
rect 833 16079 1018 16113
rect 595 16071 1018 16079
rect 595 16037 624 16071
rect 658 16041 1018 16071
rect 658 16037 799 16041
rect 595 16007 799 16037
rect 833 16007 1018 16041
rect 595 16003 1018 16007
rect 595 15969 624 16003
rect 658 15969 1018 16003
rect 595 15935 799 15969
rect 833 15935 1018 15969
rect 595 15901 624 15935
rect 658 15901 1018 15935
rect 595 15897 1018 15901
rect 595 15867 799 15897
rect 595 15833 624 15867
rect 658 15863 799 15867
rect 833 15863 1018 15897
rect 658 15833 1018 15863
rect 595 15825 1018 15833
rect 595 15799 799 15825
rect 595 15765 624 15799
rect 658 15791 799 15799
rect 833 15791 1018 15825
rect 658 15765 1018 15791
rect 595 15753 1018 15765
rect 595 15731 799 15753
rect 595 15697 624 15731
rect 658 15719 799 15731
rect 833 15719 1018 15753
rect 658 15697 1018 15719
rect 595 15681 1018 15697
rect 595 15663 799 15681
rect 595 15629 624 15663
rect 658 15647 799 15663
rect 833 15647 1018 15681
rect 658 15629 1018 15647
rect 595 15609 1018 15629
rect 595 15595 799 15609
rect 595 15561 624 15595
rect 658 15575 799 15595
rect 833 15575 1018 15609
rect 658 15561 1018 15575
rect 595 15537 1018 15561
rect 595 15527 799 15537
rect 595 15493 624 15527
rect 658 15503 799 15527
rect 833 15503 1018 15537
rect 658 15493 1018 15503
rect 595 15465 1018 15493
rect 595 15459 799 15465
rect 595 15425 624 15459
rect 658 15431 799 15459
rect 833 15431 1018 15465
rect 658 15425 1018 15431
rect 595 15393 1018 15425
rect 595 15391 799 15393
rect 595 15357 624 15391
rect 658 15359 799 15391
rect 833 15359 1018 15393
rect 658 15357 1018 15359
rect 595 15323 1018 15357
rect 595 15289 624 15323
rect 658 15321 1018 15323
rect 658 15289 799 15321
rect 595 15287 799 15289
rect 833 15287 1018 15321
rect 595 15255 1018 15287
rect 595 15221 624 15255
rect 658 15249 1018 15255
rect 658 15221 799 15249
rect 595 15215 799 15221
rect 833 15215 1018 15249
rect 595 15187 1018 15215
rect 1111 34692 13879 34734
rect 1111 34658 1293 34692
rect 1331 34658 1365 34692
rect 1399 34658 1433 34692
rect 1471 34658 1501 34692
rect 1543 34658 1569 34692
rect 1615 34658 1637 34692
rect 1687 34658 1705 34692
rect 1759 34658 1773 34692
rect 1831 34658 1841 34692
rect 1903 34658 1909 34692
rect 1975 34658 1977 34692
rect 2011 34658 2013 34692
rect 2079 34658 2085 34692
rect 2147 34658 2157 34692
rect 2215 34658 2229 34692
rect 2283 34658 2301 34692
rect 2351 34658 2373 34692
rect 2419 34658 2445 34692
rect 2487 34658 2517 34692
rect 2555 34658 2589 34692
rect 2623 34658 2657 34692
rect 2695 34658 2725 34692
rect 2767 34658 2793 34692
rect 2839 34658 2861 34692
rect 2911 34658 2929 34692
rect 2983 34658 2997 34692
rect 3055 34658 3065 34692
rect 3127 34658 3133 34692
rect 3199 34658 3201 34692
rect 3235 34658 3237 34692
rect 3303 34658 3309 34692
rect 3371 34658 3381 34692
rect 3439 34658 3453 34692
rect 3507 34658 3525 34692
rect 3575 34658 3597 34692
rect 3643 34658 3669 34692
rect 3711 34658 3741 34692
rect 3779 34658 3813 34692
rect 3847 34658 3881 34692
rect 3919 34658 3949 34692
rect 3991 34658 4017 34692
rect 4063 34658 4085 34692
rect 4135 34658 4153 34692
rect 4207 34658 4221 34692
rect 4279 34658 4289 34692
rect 4351 34658 4357 34692
rect 4423 34658 4425 34692
rect 4459 34658 4461 34692
rect 4527 34658 4533 34692
rect 4595 34658 4605 34692
rect 4663 34658 4677 34692
rect 4731 34658 4749 34692
rect 4799 34658 4821 34692
rect 4867 34658 4893 34692
rect 4935 34658 4965 34692
rect 5003 34658 5037 34692
rect 5071 34658 5105 34692
rect 5143 34658 5173 34692
rect 5215 34658 5241 34692
rect 5287 34658 5309 34692
rect 5359 34658 5377 34692
rect 5431 34658 5445 34692
rect 5503 34658 5513 34692
rect 5575 34658 5581 34692
rect 5647 34658 5649 34692
rect 5683 34658 5685 34692
rect 5751 34658 5757 34692
rect 5819 34658 5829 34692
rect 5887 34658 5901 34692
rect 5955 34658 5973 34692
rect 6023 34658 6045 34692
rect 6091 34658 6117 34692
rect 6159 34658 6189 34692
rect 6227 34658 6261 34692
rect 6295 34658 6329 34692
rect 6367 34658 6397 34692
rect 6439 34658 6465 34692
rect 6511 34658 6533 34692
rect 6583 34658 6601 34692
rect 6655 34658 6669 34692
rect 6727 34658 6737 34692
rect 6799 34658 6805 34692
rect 6871 34658 6873 34692
rect 6907 34658 6909 34692
rect 6975 34658 6981 34692
rect 7043 34658 7053 34692
rect 7111 34658 7125 34692
rect 7179 34658 7197 34692
rect 7247 34658 7269 34692
rect 7315 34658 7341 34692
rect 7383 34658 7413 34692
rect 7451 34658 7485 34692
rect 7519 34658 7553 34692
rect 7591 34658 7621 34692
rect 7663 34658 7689 34692
rect 7735 34658 7757 34692
rect 7807 34658 7825 34692
rect 7879 34658 7893 34692
rect 7951 34658 7961 34692
rect 8023 34658 8029 34692
rect 8095 34658 8097 34692
rect 8131 34658 8133 34692
rect 8199 34658 8205 34692
rect 8267 34658 8277 34692
rect 8335 34658 8349 34692
rect 8403 34658 8421 34692
rect 8471 34658 8493 34692
rect 8539 34658 8565 34692
rect 8607 34658 8637 34692
rect 8675 34658 8709 34692
rect 8743 34658 8777 34692
rect 8815 34658 8845 34692
rect 8887 34658 8913 34692
rect 8959 34658 8981 34692
rect 9031 34658 9049 34692
rect 9103 34658 9117 34692
rect 9175 34658 9185 34692
rect 9247 34658 9253 34692
rect 9319 34658 9321 34692
rect 9355 34658 9357 34692
rect 9423 34658 9429 34692
rect 9491 34658 9501 34692
rect 9559 34658 9573 34692
rect 9627 34658 9645 34692
rect 9695 34658 9717 34692
rect 9763 34658 9789 34692
rect 9831 34658 9861 34692
rect 9899 34658 9933 34692
rect 9967 34658 10001 34692
rect 10039 34658 10069 34692
rect 10111 34658 10137 34692
rect 10183 34658 10205 34692
rect 10255 34658 10273 34692
rect 10327 34658 10341 34692
rect 10399 34658 10409 34692
rect 10471 34658 10477 34692
rect 10543 34658 10545 34692
rect 10579 34658 10581 34692
rect 10647 34658 10653 34692
rect 10715 34658 10725 34692
rect 10783 34658 10797 34692
rect 10851 34658 10869 34692
rect 10919 34658 10941 34692
rect 10987 34658 11013 34692
rect 11055 34658 11085 34692
rect 11123 34658 11157 34692
rect 11191 34658 11225 34692
rect 11263 34658 11293 34692
rect 11335 34658 11361 34692
rect 11407 34658 11429 34692
rect 11479 34658 11497 34692
rect 11551 34658 11565 34692
rect 11623 34658 11633 34692
rect 11695 34658 11701 34692
rect 11767 34658 11769 34692
rect 11803 34658 11805 34692
rect 11871 34658 11877 34692
rect 11939 34658 11949 34692
rect 12007 34658 12021 34692
rect 12075 34658 12093 34692
rect 12143 34658 12165 34692
rect 12211 34658 12237 34692
rect 12279 34658 12309 34692
rect 12347 34658 12381 34692
rect 12415 34658 12449 34692
rect 12487 34658 12517 34692
rect 12559 34658 12585 34692
rect 12631 34658 12653 34692
rect 12703 34658 12721 34692
rect 12775 34658 12789 34692
rect 12847 34658 12857 34692
rect 12919 34658 12925 34692
rect 12991 34658 12993 34692
rect 13027 34658 13029 34692
rect 13095 34658 13101 34692
rect 13163 34658 13173 34692
rect 13231 34658 13245 34692
rect 13299 34658 13317 34692
rect 13367 34658 13389 34692
rect 13435 34658 13461 34692
rect 13503 34658 13533 34692
rect 13571 34658 13605 34692
rect 13639 34658 13673 34692
rect 13711 34658 13879 34692
rect 1111 34616 13879 34658
rect 1111 34495 1229 34616
rect 1111 34441 1153 34495
rect 1187 34441 1229 34495
rect 1111 34423 1229 34441
rect 1111 34373 1153 34423
rect 1187 34373 1229 34423
rect 1111 34351 1229 34373
rect 1111 34305 1153 34351
rect 1187 34305 1229 34351
rect 1111 34279 1229 34305
rect 1111 34237 1153 34279
rect 1187 34237 1229 34279
rect 1111 34207 1229 34237
rect 1111 34169 1153 34207
rect 1187 34169 1229 34207
rect 1111 34135 1229 34169
rect 1111 34101 1153 34135
rect 1187 34101 1229 34135
rect 1111 34067 1229 34101
rect 1111 34029 1153 34067
rect 1187 34029 1229 34067
rect 1111 33999 1229 34029
rect 1111 33957 1153 33999
rect 1187 33957 1229 33999
rect 1111 33931 1229 33957
rect 1111 33885 1153 33931
rect 1187 33885 1229 33931
rect 1111 33863 1229 33885
rect 1111 33813 1153 33863
rect 1187 33813 1229 33863
rect 1111 33795 1229 33813
rect 1111 33741 1153 33795
rect 1187 33741 1229 33795
rect 1111 33727 1229 33741
rect 1111 33669 1153 33727
rect 1187 33669 1229 33727
rect 1111 33659 1229 33669
rect 1111 33597 1153 33659
rect 1187 33597 1229 33659
rect 1111 33591 1229 33597
rect 1111 33525 1153 33591
rect 1187 33525 1229 33591
rect 1111 33523 1229 33525
rect 1111 33489 1153 33523
rect 1187 33489 1229 33523
rect 1111 33487 1229 33489
rect 1111 33421 1153 33487
rect 1187 33421 1229 33487
rect 1111 33415 1229 33421
rect 1111 33353 1153 33415
rect 1187 33353 1229 33415
rect 1111 33343 1229 33353
rect 1111 33285 1153 33343
rect 1187 33285 1229 33343
rect 1111 33271 1229 33285
rect 1111 33217 1153 33271
rect 1187 33217 1229 33271
rect 1111 33199 1229 33217
rect 1111 33149 1153 33199
rect 1187 33149 1229 33199
rect 1111 33127 1229 33149
rect 1111 33081 1153 33127
rect 1187 33081 1229 33127
rect 1111 33055 1229 33081
rect 1111 33013 1153 33055
rect 1187 33013 1229 33055
rect 1111 32983 1229 33013
rect 1111 32945 1153 32983
rect 1187 32945 1229 32983
rect 1111 32911 1229 32945
rect 1111 32877 1153 32911
rect 1187 32877 1229 32911
rect 1111 32843 1229 32877
rect 1111 32805 1153 32843
rect 1187 32805 1229 32843
rect 1111 32775 1229 32805
rect 1111 32733 1153 32775
rect 1187 32733 1229 32775
rect 1111 32707 1229 32733
rect 1111 32661 1153 32707
rect 1187 32661 1229 32707
rect 1111 32639 1229 32661
rect 1111 32589 1153 32639
rect 1187 32589 1229 32639
rect 1111 32571 1229 32589
rect 1111 32517 1153 32571
rect 1187 32517 1229 32571
rect 1111 32503 1229 32517
rect 1111 32445 1153 32503
rect 1187 32445 1229 32503
rect 1111 32435 1229 32445
rect 1111 32373 1153 32435
rect 1187 32373 1229 32435
rect 1111 32367 1229 32373
rect 1111 32301 1153 32367
rect 1187 32301 1229 32367
rect 1111 32299 1229 32301
rect 1111 32265 1153 32299
rect 1187 32265 1229 32299
rect 1111 32263 1229 32265
rect 1111 32197 1153 32263
rect 1187 32197 1229 32263
rect 1111 32191 1229 32197
rect 1111 32129 1153 32191
rect 1187 32129 1229 32191
rect 1111 32119 1229 32129
rect 1111 32061 1153 32119
rect 1187 32061 1229 32119
rect 1111 32047 1229 32061
rect 1111 31993 1153 32047
rect 1187 31993 1229 32047
rect 1111 31975 1229 31993
rect 1111 31925 1153 31975
rect 1187 31925 1229 31975
rect 1111 31903 1229 31925
rect 1111 31857 1153 31903
rect 1187 31857 1229 31903
rect 1111 31831 1229 31857
rect 1111 31789 1153 31831
rect 1187 31789 1229 31831
rect 1111 31759 1229 31789
rect 1111 31721 1153 31759
rect 1187 31721 1229 31759
rect 1111 31687 1229 31721
rect 1111 31653 1153 31687
rect 1187 31653 1229 31687
rect 1111 31619 1229 31653
rect 1111 31581 1153 31619
rect 1187 31581 1229 31619
rect 1111 31551 1229 31581
rect 1111 31509 1153 31551
rect 1187 31509 1229 31551
rect 1111 31483 1229 31509
rect 1111 31437 1153 31483
rect 1187 31437 1229 31483
rect 1111 31415 1229 31437
rect 1111 31365 1153 31415
rect 1187 31365 1229 31415
rect 1111 31347 1229 31365
rect 1111 31293 1153 31347
rect 1187 31293 1229 31347
rect 1111 31279 1229 31293
rect 1111 31221 1153 31279
rect 1187 31221 1229 31279
rect 1111 31211 1229 31221
rect 1111 31149 1153 31211
rect 1187 31149 1229 31211
rect 1111 31143 1229 31149
rect 1111 31077 1153 31143
rect 1187 31077 1229 31143
rect 1111 31075 1229 31077
rect 1111 31041 1153 31075
rect 1187 31041 1229 31075
rect 1111 31039 1229 31041
rect 1111 30973 1153 31039
rect 1187 30973 1229 31039
rect 1111 30967 1229 30973
rect 1111 30905 1153 30967
rect 1187 30905 1229 30967
rect 1111 30895 1229 30905
rect 1111 30837 1153 30895
rect 1187 30837 1229 30895
rect 1111 30823 1229 30837
rect 1111 30769 1153 30823
rect 1187 30769 1229 30823
rect 1111 30751 1229 30769
rect 1111 30701 1153 30751
rect 1187 30701 1229 30751
rect 1111 30679 1229 30701
rect 1111 30633 1153 30679
rect 1187 30633 1229 30679
rect 1111 30607 1229 30633
rect 1111 30565 1153 30607
rect 1187 30565 1229 30607
rect 1111 30535 1229 30565
rect 1111 30497 1153 30535
rect 1187 30497 1229 30535
rect 1111 30463 1229 30497
rect 1111 30429 1153 30463
rect 1187 30429 1229 30463
rect 1111 30395 1229 30429
rect 1111 30357 1153 30395
rect 1187 30357 1229 30395
rect 1111 30327 1229 30357
rect 1111 30285 1153 30327
rect 1187 30285 1229 30327
rect 1111 30259 1229 30285
rect 1111 30213 1153 30259
rect 1187 30213 1229 30259
rect 1111 30191 1229 30213
rect 1111 30141 1153 30191
rect 1187 30141 1229 30191
rect 1111 30123 1229 30141
rect 1111 30069 1153 30123
rect 1187 30069 1229 30123
rect 1111 30055 1229 30069
rect 1111 29997 1153 30055
rect 1187 29997 1229 30055
rect 1111 29987 1229 29997
rect 1111 29925 1153 29987
rect 1187 29925 1229 29987
rect 1111 29919 1229 29925
rect 1111 29853 1153 29919
rect 1187 29853 1229 29919
rect 1111 29851 1229 29853
rect 1111 29817 1153 29851
rect 1187 29817 1229 29851
rect 1111 29815 1229 29817
rect 1111 29749 1153 29815
rect 1187 29749 1229 29815
rect 1111 29743 1229 29749
rect 1111 29681 1153 29743
rect 1187 29681 1229 29743
rect 1111 29671 1229 29681
rect 1111 29613 1153 29671
rect 1187 29613 1229 29671
rect 1111 29599 1229 29613
rect 1111 29545 1153 29599
rect 1187 29545 1229 29599
rect 1111 29527 1229 29545
rect 1111 29477 1153 29527
rect 1187 29477 1229 29527
rect 1111 29455 1229 29477
rect 1111 29409 1153 29455
rect 1187 29409 1229 29455
rect 1111 29383 1229 29409
rect 1111 29341 1153 29383
rect 1187 29341 1229 29383
rect 1111 29311 1229 29341
rect 1111 29273 1153 29311
rect 1187 29273 1229 29311
rect 1111 29239 1229 29273
rect 1111 29205 1153 29239
rect 1187 29205 1229 29239
rect 1111 29171 1229 29205
rect 1111 29133 1153 29171
rect 1187 29133 1229 29171
rect 1111 29103 1229 29133
rect 1111 29061 1153 29103
rect 1187 29061 1229 29103
rect 1111 29035 1229 29061
rect 1111 28989 1153 29035
rect 1187 28989 1229 29035
rect 1111 28967 1229 28989
rect 1111 28917 1153 28967
rect 1187 28917 1229 28967
rect 13761 34487 13879 34616
rect 13761 34436 13801 34487
rect 13835 34436 13879 34487
rect 13761 34415 13879 34436
rect 13761 34368 13801 34415
rect 13835 34368 13879 34415
rect 13761 34343 13879 34368
rect 13761 34300 13801 34343
rect 13835 34300 13879 34343
rect 13761 34271 13879 34300
rect 13761 34232 13801 34271
rect 13835 34232 13879 34271
rect 13761 34199 13879 34232
rect 13761 34164 13801 34199
rect 13835 34164 13879 34199
rect 13761 34130 13879 34164
rect 13761 34093 13801 34130
rect 13835 34093 13879 34130
rect 13761 34062 13879 34093
rect 13761 34021 13801 34062
rect 13835 34021 13879 34062
rect 13761 33994 13879 34021
rect 13761 33949 13801 33994
rect 13835 33949 13879 33994
rect 13761 33926 13879 33949
rect 13761 33877 13801 33926
rect 13835 33877 13879 33926
rect 13761 33858 13879 33877
rect 13761 33805 13801 33858
rect 13835 33805 13879 33858
rect 13761 33790 13879 33805
rect 13761 33733 13801 33790
rect 13835 33733 13879 33790
rect 13761 33722 13879 33733
rect 13761 33661 13801 33722
rect 13835 33661 13879 33722
rect 13761 33654 13879 33661
rect 13761 33589 13801 33654
rect 13835 33589 13879 33654
rect 13761 33586 13879 33589
rect 13761 33552 13801 33586
rect 13835 33552 13879 33586
rect 13761 33551 13879 33552
rect 13761 33484 13801 33551
rect 13835 33484 13879 33551
rect 13761 33479 13879 33484
rect 13761 33416 13801 33479
rect 13835 33416 13879 33479
rect 13761 33407 13879 33416
rect 13761 33348 13801 33407
rect 13835 33348 13879 33407
rect 13761 33335 13879 33348
rect 13761 33280 13801 33335
rect 13835 33280 13879 33335
rect 13761 33263 13879 33280
rect 13761 33212 13801 33263
rect 13835 33212 13879 33263
rect 13761 33191 13879 33212
rect 13761 33144 13801 33191
rect 13835 33144 13879 33191
rect 13761 33119 13879 33144
rect 13761 33076 13801 33119
rect 13835 33076 13879 33119
rect 13761 33047 13879 33076
rect 13761 33008 13801 33047
rect 13835 33008 13879 33047
rect 13761 32975 13879 33008
rect 13761 32940 13801 32975
rect 13835 32940 13879 32975
rect 13761 32906 13879 32940
rect 13761 32869 13801 32906
rect 13835 32869 13879 32906
rect 13761 32838 13879 32869
rect 13761 32797 13801 32838
rect 13835 32797 13879 32838
rect 13761 32770 13879 32797
rect 13761 32725 13801 32770
rect 13835 32725 13879 32770
rect 13761 32702 13879 32725
rect 13761 32653 13801 32702
rect 13835 32653 13879 32702
rect 13761 32634 13879 32653
rect 13761 32581 13801 32634
rect 13835 32581 13879 32634
rect 13761 32566 13879 32581
rect 13761 32509 13801 32566
rect 13835 32509 13879 32566
rect 13761 32498 13879 32509
rect 13761 32437 13801 32498
rect 13835 32437 13879 32498
rect 13761 32430 13879 32437
rect 13761 32365 13801 32430
rect 13835 32365 13879 32430
rect 13761 32362 13879 32365
rect 13761 32328 13801 32362
rect 13835 32328 13879 32362
rect 13761 32327 13879 32328
rect 13761 32260 13801 32327
rect 13835 32260 13879 32327
rect 13761 32255 13879 32260
rect 13761 32192 13801 32255
rect 13835 32192 13879 32255
rect 13761 32183 13879 32192
rect 13761 32124 13801 32183
rect 13835 32124 13879 32183
rect 13761 32111 13879 32124
rect 13761 32056 13801 32111
rect 13835 32056 13879 32111
rect 13761 32039 13879 32056
rect 13761 31988 13801 32039
rect 13835 31988 13879 32039
rect 13761 31967 13879 31988
rect 13761 31920 13801 31967
rect 13835 31920 13879 31967
rect 13761 31895 13879 31920
rect 13761 31852 13801 31895
rect 13835 31852 13879 31895
rect 13761 31823 13879 31852
rect 13761 31784 13801 31823
rect 13835 31784 13879 31823
rect 13761 31751 13879 31784
rect 13761 31716 13801 31751
rect 13835 31716 13879 31751
rect 13761 31682 13879 31716
rect 13761 31645 13801 31682
rect 13835 31645 13879 31682
rect 13761 31614 13879 31645
rect 13761 31573 13801 31614
rect 13835 31573 13879 31614
rect 13761 31546 13879 31573
rect 13761 31501 13801 31546
rect 13835 31501 13879 31546
rect 13761 31478 13879 31501
rect 13761 31429 13801 31478
rect 13835 31429 13879 31478
rect 13761 31410 13879 31429
rect 13761 31357 13801 31410
rect 13835 31357 13879 31410
rect 13761 31342 13879 31357
rect 13761 31285 13801 31342
rect 13835 31285 13879 31342
rect 13761 31274 13879 31285
rect 13761 31213 13801 31274
rect 13835 31213 13879 31274
rect 13761 31206 13879 31213
rect 13761 31141 13801 31206
rect 13835 31141 13879 31206
rect 13761 31138 13879 31141
rect 13761 31104 13801 31138
rect 13835 31104 13879 31138
rect 13761 31103 13879 31104
rect 13761 31036 13801 31103
rect 13835 31036 13879 31103
rect 13761 31031 13879 31036
rect 13761 30968 13801 31031
rect 13835 30968 13879 31031
rect 13761 30959 13879 30968
rect 13761 30900 13801 30959
rect 13835 30900 13879 30959
rect 13761 30887 13879 30900
rect 13761 30832 13801 30887
rect 13835 30832 13879 30887
rect 13761 30815 13879 30832
rect 13761 30764 13801 30815
rect 13835 30764 13879 30815
rect 13761 30743 13879 30764
rect 13761 30696 13801 30743
rect 13835 30696 13879 30743
rect 13761 30671 13879 30696
rect 13761 30628 13801 30671
rect 13835 30628 13879 30671
rect 13761 30599 13879 30628
rect 13761 30560 13801 30599
rect 13835 30560 13879 30599
rect 13761 30527 13879 30560
rect 13761 30492 13801 30527
rect 13835 30492 13879 30527
rect 13761 30458 13879 30492
rect 13761 30421 13801 30458
rect 13835 30421 13879 30458
rect 13761 30390 13879 30421
rect 13761 30349 13801 30390
rect 13835 30349 13879 30390
rect 13761 30322 13879 30349
rect 13761 30277 13801 30322
rect 13835 30277 13879 30322
rect 13761 30254 13879 30277
rect 13761 30205 13801 30254
rect 13835 30205 13879 30254
rect 13761 30186 13879 30205
rect 13761 30133 13801 30186
rect 13835 30133 13879 30186
rect 13761 30118 13879 30133
rect 13761 30061 13801 30118
rect 13835 30061 13879 30118
rect 13761 30050 13879 30061
rect 13761 29989 13801 30050
rect 13835 29989 13879 30050
rect 13761 29982 13879 29989
rect 13761 29917 13801 29982
rect 13835 29917 13879 29982
rect 13761 29914 13879 29917
rect 13761 29880 13801 29914
rect 13835 29880 13879 29914
rect 13761 29879 13879 29880
rect 13761 29812 13801 29879
rect 13835 29812 13879 29879
rect 13761 29807 13879 29812
rect 13761 29744 13801 29807
rect 13835 29744 13879 29807
rect 13761 29735 13879 29744
rect 13761 29676 13801 29735
rect 13835 29676 13879 29735
rect 13761 29663 13879 29676
rect 13761 29608 13801 29663
rect 13835 29608 13879 29663
rect 13761 29591 13879 29608
rect 13761 29540 13801 29591
rect 13835 29540 13879 29591
rect 13761 29519 13879 29540
rect 13761 29472 13801 29519
rect 13835 29472 13879 29519
rect 13761 29447 13879 29472
rect 13761 29404 13801 29447
rect 13835 29404 13879 29447
rect 13761 29375 13879 29404
rect 13761 29336 13801 29375
rect 13835 29336 13879 29375
rect 13761 29303 13879 29336
rect 13761 29268 13801 29303
rect 13835 29268 13879 29303
rect 13761 29234 13879 29268
rect 13761 29197 13801 29234
rect 13835 29197 13879 29234
rect 13761 29166 13879 29197
rect 13761 29125 13801 29166
rect 13835 29125 13879 29166
rect 13761 29098 13879 29125
rect 13761 29053 13801 29098
rect 13835 29053 13879 29098
rect 13761 29030 13879 29053
rect 13761 28981 13801 29030
rect 13835 28981 13879 29030
rect 13761 28962 13879 28981
rect 1111 28899 1229 28917
rect 1111 28845 1153 28899
rect 1187 28845 1229 28899
rect 1111 28831 1229 28845
rect 1111 28773 1153 28831
rect 1187 28773 1229 28831
rect 1111 28763 1229 28773
rect 1111 28701 1153 28763
rect 1187 28701 1229 28763
rect 1111 28695 1229 28701
rect 1111 28629 1153 28695
rect 1187 28629 1229 28695
rect 1111 28627 1229 28629
rect 1111 28593 1153 28627
rect 1187 28593 1229 28627
rect 1111 28591 1229 28593
rect 1111 28525 1153 28591
rect 1187 28525 1229 28591
rect 1111 28519 1229 28525
rect 1111 28457 1153 28519
rect 1187 28457 1229 28519
rect 1111 28447 1229 28457
rect 1111 28389 1153 28447
rect 1187 28389 1229 28447
rect 1111 28375 1229 28389
rect 1111 28321 1153 28375
rect 1187 28321 1229 28375
rect 1111 28303 1229 28321
rect 1111 28253 1153 28303
rect 1187 28253 1229 28303
rect 1111 28231 1229 28253
rect 1111 28185 1153 28231
rect 1187 28185 1229 28231
rect 1111 28159 1229 28185
rect 1111 28117 1153 28159
rect 1187 28117 1229 28159
rect 1111 28087 1229 28117
rect 1111 28049 1153 28087
rect 1187 28049 1229 28087
rect 1111 28015 1229 28049
rect 1111 27981 1153 28015
rect 1187 27981 1229 28015
rect 1111 27947 1229 27981
rect 1111 27909 1153 27947
rect 1187 27909 1229 27947
rect 1111 27879 1229 27909
rect 1111 27837 1153 27879
rect 1187 27837 1229 27879
rect 1111 27811 1229 27837
rect 1111 27765 1153 27811
rect 1187 27765 1229 27811
rect 1111 27743 1229 27765
rect 1111 27693 1153 27743
rect 1187 27693 1229 27743
rect 1111 27675 1229 27693
rect 1111 27621 1153 27675
rect 1187 27621 1229 27675
rect 1111 27607 1229 27621
rect 1111 27549 1153 27607
rect 1187 27549 1229 27607
rect 1111 27539 1229 27549
rect 1111 27477 1153 27539
rect 1187 27477 1229 27539
rect 1111 27471 1229 27477
rect 1111 27405 1153 27471
rect 1187 27405 1229 27471
rect 1111 27403 1229 27405
rect 1111 27369 1153 27403
rect 1187 27369 1229 27403
rect 1111 27367 1229 27369
rect 1111 27301 1153 27367
rect 1187 27301 1229 27367
rect 1111 27295 1229 27301
rect 1111 27233 1153 27295
rect 1187 27233 1229 27295
rect 1111 27223 1229 27233
rect 1111 27165 1153 27223
rect 1187 27165 1229 27223
rect 1111 27151 1229 27165
rect 1111 27097 1153 27151
rect 1187 27097 1229 27151
rect 1111 27079 1229 27097
rect 1111 27029 1153 27079
rect 1187 27029 1229 27079
rect 1651 28892 13349 28922
rect 1651 28888 2111 28892
rect 12889 28888 13349 28892
rect 1651 28566 1974 28888
rect 13024 28566 13349 28888
rect 1651 28518 2111 28566
rect 12889 28518 13349 28566
rect 1651 28502 13349 28518
rect 1651 28435 1718 28502
rect 1968 28495 13349 28502
rect 1968 28488 13023 28495
rect 1968 28435 2085 28488
rect 1651 27517 1681 28435
rect 2055 27517 2085 28435
rect 12915 28435 13023 28488
rect 13273 28435 13349 28495
rect 2148 28277 12832 28381
rect 2148 28243 2443 28277
rect 2477 28273 2515 28277
rect 2549 28273 2587 28277
rect 2477 28243 2485 28273
rect 2549 28243 2553 28273
rect 2148 28239 2485 28243
rect 2519 28239 2553 28243
rect 2621 28273 2659 28277
rect 2693 28273 2731 28277
rect 2765 28273 2803 28277
rect 2837 28273 2875 28277
rect 2909 28273 2947 28277
rect 2981 28273 3019 28277
rect 3053 28273 3091 28277
rect 3125 28273 3163 28277
rect 3197 28273 3235 28277
rect 3269 28273 3307 28277
rect 3341 28273 3379 28277
rect 3413 28273 3451 28277
rect 3485 28273 3523 28277
rect 3557 28273 3595 28277
rect 3629 28273 3667 28277
rect 3701 28273 3739 28277
rect 3773 28273 3811 28277
rect 2587 28239 2621 28243
rect 2655 28243 2659 28273
rect 2723 28243 2731 28273
rect 2791 28243 2803 28273
rect 2859 28243 2875 28273
rect 2927 28243 2947 28273
rect 2995 28243 3019 28273
rect 3063 28243 3091 28273
rect 3131 28243 3163 28273
rect 2655 28239 2689 28243
rect 2723 28239 2757 28243
rect 2791 28239 2825 28243
rect 2859 28239 2893 28243
rect 2927 28239 2961 28243
rect 2995 28239 3029 28243
rect 3063 28239 3097 28243
rect 3131 28239 3165 28243
rect 3199 28239 3233 28273
rect 3269 28243 3301 28273
rect 3341 28243 3369 28273
rect 3413 28243 3437 28273
rect 3485 28243 3505 28273
rect 3557 28243 3573 28273
rect 3629 28243 3641 28273
rect 3701 28243 3709 28273
rect 3773 28243 3777 28273
rect 3267 28239 3301 28243
rect 3335 28239 3369 28243
rect 3403 28239 3437 28243
rect 3471 28239 3505 28243
rect 3539 28239 3573 28243
rect 3607 28239 3641 28243
rect 3675 28239 3709 28243
rect 3743 28239 3777 28243
rect 3845 28273 3883 28277
rect 3917 28273 3955 28277
rect 3989 28273 4027 28277
rect 4061 28273 4099 28277
rect 4133 28273 4171 28277
rect 4205 28273 4243 28277
rect 4277 28273 4315 28277
rect 4349 28273 4387 28277
rect 4421 28273 4459 28277
rect 4493 28273 4531 28277
rect 4565 28273 4603 28277
rect 4637 28273 4675 28277
rect 4709 28273 4747 28277
rect 4781 28273 4819 28277
rect 4853 28273 4891 28277
rect 4925 28273 4963 28277
rect 4997 28273 5035 28277
rect 3811 28239 3845 28243
rect 3879 28243 3883 28273
rect 3947 28243 3955 28273
rect 4015 28243 4027 28273
rect 4083 28243 4099 28273
rect 4151 28243 4171 28273
rect 4219 28243 4243 28273
rect 4287 28243 4315 28273
rect 4355 28243 4387 28273
rect 3879 28239 3913 28243
rect 3947 28239 3981 28243
rect 4015 28239 4049 28243
rect 4083 28239 4117 28243
rect 4151 28239 4185 28243
rect 4219 28239 4253 28243
rect 4287 28239 4321 28243
rect 4355 28239 4389 28243
rect 4423 28239 4457 28273
rect 4493 28243 4525 28273
rect 4565 28243 4593 28273
rect 4637 28243 4661 28273
rect 4709 28243 4729 28273
rect 4781 28243 4797 28273
rect 4853 28243 4865 28273
rect 4925 28243 4933 28273
rect 4997 28243 5001 28273
rect 4491 28239 4525 28243
rect 4559 28239 4593 28243
rect 4627 28239 4661 28243
rect 4695 28239 4729 28243
rect 4763 28239 4797 28243
rect 4831 28239 4865 28243
rect 4899 28239 4933 28243
rect 4967 28239 5001 28243
rect 5069 28273 5107 28277
rect 5141 28273 5179 28277
rect 5213 28273 5251 28277
rect 5285 28273 5323 28277
rect 5357 28273 5395 28277
rect 5429 28273 5467 28277
rect 5501 28273 5539 28277
rect 5573 28273 5611 28277
rect 5645 28273 5683 28277
rect 5717 28273 5755 28277
rect 5789 28273 5827 28277
rect 5861 28273 5899 28277
rect 5933 28273 5971 28277
rect 6005 28273 6043 28277
rect 6077 28273 6115 28277
rect 6149 28273 6187 28277
rect 6221 28273 6259 28277
rect 5035 28239 5069 28243
rect 5103 28243 5107 28273
rect 5171 28243 5179 28273
rect 5239 28243 5251 28273
rect 5307 28243 5323 28273
rect 5375 28243 5395 28273
rect 5443 28243 5467 28273
rect 5511 28243 5539 28273
rect 5579 28243 5611 28273
rect 5103 28239 5137 28243
rect 5171 28239 5205 28243
rect 5239 28239 5273 28243
rect 5307 28239 5341 28243
rect 5375 28239 5409 28243
rect 5443 28239 5477 28243
rect 5511 28239 5545 28243
rect 5579 28239 5613 28243
rect 5647 28239 5681 28273
rect 5717 28243 5749 28273
rect 5789 28243 5817 28273
rect 5861 28243 5885 28273
rect 5933 28243 5953 28273
rect 6005 28243 6021 28273
rect 6077 28243 6089 28273
rect 6149 28243 6157 28273
rect 6221 28243 6225 28273
rect 5715 28239 5749 28243
rect 5783 28239 5817 28243
rect 5851 28239 5885 28243
rect 5919 28239 5953 28243
rect 5987 28239 6021 28243
rect 6055 28239 6089 28243
rect 6123 28239 6157 28243
rect 6191 28239 6225 28243
rect 6293 28273 6331 28277
rect 6365 28273 6403 28277
rect 6437 28273 6475 28277
rect 6509 28273 6547 28277
rect 6581 28273 6619 28277
rect 6653 28273 6691 28277
rect 6725 28273 6763 28277
rect 6797 28273 6835 28277
rect 6869 28273 6907 28277
rect 6941 28273 6979 28277
rect 7013 28273 7051 28277
rect 7085 28273 7123 28277
rect 7157 28273 7195 28277
rect 7229 28273 7267 28277
rect 7301 28273 7339 28277
rect 7373 28273 7411 28277
rect 7445 28273 7483 28277
rect 6259 28239 6293 28243
rect 6327 28243 6331 28273
rect 6395 28243 6403 28273
rect 6463 28243 6475 28273
rect 6531 28243 6547 28273
rect 6599 28243 6619 28273
rect 6667 28243 6691 28273
rect 6735 28243 6763 28273
rect 6803 28243 6835 28273
rect 6327 28239 6361 28243
rect 6395 28239 6429 28243
rect 6463 28239 6497 28243
rect 6531 28239 6565 28243
rect 6599 28239 6633 28243
rect 6667 28239 6701 28243
rect 6735 28239 6769 28243
rect 6803 28239 6837 28243
rect 6871 28239 6905 28273
rect 6941 28243 6973 28273
rect 7013 28243 7041 28273
rect 7085 28243 7109 28273
rect 7157 28243 7177 28273
rect 7229 28243 7245 28273
rect 7301 28243 7313 28273
rect 7373 28243 7381 28273
rect 7445 28243 7449 28273
rect 6939 28239 6973 28243
rect 7007 28239 7041 28243
rect 7075 28239 7109 28243
rect 7143 28239 7177 28243
rect 7211 28239 7245 28243
rect 7279 28239 7313 28243
rect 7347 28239 7381 28243
rect 7415 28239 7449 28243
rect 7517 28273 7555 28277
rect 7589 28273 7627 28277
rect 7661 28273 7699 28277
rect 7733 28273 7771 28277
rect 7805 28273 7843 28277
rect 7877 28273 7915 28277
rect 7949 28273 7987 28277
rect 8021 28273 8059 28277
rect 8093 28273 8131 28277
rect 8165 28273 8203 28277
rect 8237 28273 8275 28277
rect 8309 28273 8347 28277
rect 8381 28273 8419 28277
rect 8453 28273 8491 28277
rect 8525 28273 8563 28277
rect 8597 28273 8635 28277
rect 8669 28273 8707 28277
rect 7483 28239 7517 28243
rect 7551 28243 7555 28273
rect 7619 28243 7627 28273
rect 7687 28243 7699 28273
rect 7755 28243 7771 28273
rect 7823 28243 7843 28273
rect 7891 28243 7915 28273
rect 7959 28243 7987 28273
rect 8027 28243 8059 28273
rect 7551 28239 7585 28243
rect 7619 28239 7653 28243
rect 7687 28239 7721 28243
rect 7755 28239 7789 28243
rect 7823 28239 7857 28243
rect 7891 28239 7925 28243
rect 7959 28239 7993 28243
rect 8027 28239 8061 28243
rect 8095 28239 8129 28273
rect 8165 28243 8197 28273
rect 8237 28243 8265 28273
rect 8309 28243 8333 28273
rect 8381 28243 8401 28273
rect 8453 28243 8469 28273
rect 8525 28243 8537 28273
rect 8597 28243 8605 28273
rect 8669 28243 8673 28273
rect 8163 28239 8197 28243
rect 8231 28239 8265 28243
rect 8299 28239 8333 28243
rect 8367 28239 8401 28243
rect 8435 28239 8469 28243
rect 8503 28239 8537 28243
rect 8571 28239 8605 28243
rect 8639 28239 8673 28243
rect 8741 28273 8779 28277
rect 8813 28273 8851 28277
rect 8885 28273 8923 28277
rect 8957 28273 8995 28277
rect 9029 28273 9067 28277
rect 9101 28273 9139 28277
rect 9173 28273 9211 28277
rect 9245 28273 9283 28277
rect 9317 28273 9355 28277
rect 9389 28273 9427 28277
rect 9461 28273 9499 28277
rect 9533 28273 9571 28277
rect 9605 28273 9643 28277
rect 9677 28273 9715 28277
rect 9749 28273 9787 28277
rect 9821 28273 9859 28277
rect 9893 28273 9931 28277
rect 8707 28239 8741 28243
rect 8775 28243 8779 28273
rect 8843 28243 8851 28273
rect 8911 28243 8923 28273
rect 8979 28243 8995 28273
rect 9047 28243 9067 28273
rect 9115 28243 9139 28273
rect 9183 28243 9211 28273
rect 9251 28243 9283 28273
rect 8775 28239 8809 28243
rect 8843 28239 8877 28243
rect 8911 28239 8945 28243
rect 8979 28239 9013 28243
rect 9047 28239 9081 28243
rect 9115 28239 9149 28243
rect 9183 28239 9217 28243
rect 9251 28239 9285 28243
rect 9319 28239 9353 28273
rect 9389 28243 9421 28273
rect 9461 28243 9489 28273
rect 9533 28243 9557 28273
rect 9605 28243 9625 28273
rect 9677 28243 9693 28273
rect 9749 28243 9761 28273
rect 9821 28243 9829 28273
rect 9893 28243 9897 28273
rect 9387 28239 9421 28243
rect 9455 28239 9489 28243
rect 9523 28239 9557 28243
rect 9591 28239 9625 28243
rect 9659 28239 9693 28243
rect 9727 28239 9761 28243
rect 9795 28239 9829 28243
rect 9863 28239 9897 28243
rect 9965 28273 10003 28277
rect 10037 28273 10075 28277
rect 10109 28273 10147 28277
rect 10181 28273 10219 28277
rect 10253 28273 10291 28277
rect 10325 28273 10363 28277
rect 10397 28273 10435 28277
rect 10469 28273 10507 28277
rect 10541 28273 10579 28277
rect 10613 28273 10651 28277
rect 10685 28273 10723 28277
rect 10757 28273 10795 28277
rect 10829 28273 10867 28277
rect 10901 28273 10939 28277
rect 10973 28273 11011 28277
rect 11045 28273 11083 28277
rect 11117 28273 11155 28277
rect 9931 28239 9965 28243
rect 9999 28243 10003 28273
rect 10067 28243 10075 28273
rect 10135 28243 10147 28273
rect 10203 28243 10219 28273
rect 10271 28243 10291 28273
rect 10339 28243 10363 28273
rect 10407 28243 10435 28273
rect 10475 28243 10507 28273
rect 9999 28239 10033 28243
rect 10067 28239 10101 28243
rect 10135 28239 10169 28243
rect 10203 28239 10237 28243
rect 10271 28239 10305 28243
rect 10339 28239 10373 28243
rect 10407 28239 10441 28243
rect 10475 28239 10509 28243
rect 10543 28239 10577 28273
rect 10613 28243 10645 28273
rect 10685 28243 10713 28273
rect 10757 28243 10781 28273
rect 10829 28243 10849 28273
rect 10901 28243 10917 28273
rect 10973 28243 10985 28273
rect 11045 28243 11053 28273
rect 11117 28243 11121 28273
rect 10611 28239 10645 28243
rect 10679 28239 10713 28243
rect 10747 28239 10781 28243
rect 10815 28239 10849 28243
rect 10883 28239 10917 28243
rect 10951 28239 10985 28243
rect 11019 28239 11053 28243
rect 11087 28239 11121 28243
rect 11189 28273 11227 28277
rect 11261 28273 11299 28277
rect 11333 28273 11371 28277
rect 11405 28273 11443 28277
rect 11477 28273 11515 28277
rect 11549 28273 11587 28277
rect 11621 28273 11659 28277
rect 11693 28273 11731 28277
rect 11765 28273 11803 28277
rect 11837 28273 11875 28277
rect 11909 28273 11947 28277
rect 11981 28273 12019 28277
rect 12053 28273 12091 28277
rect 12125 28273 12163 28277
rect 12197 28273 12235 28277
rect 12269 28273 12307 28277
rect 12341 28273 12379 28277
rect 11155 28239 11189 28243
rect 11223 28243 11227 28273
rect 11291 28243 11299 28273
rect 11359 28243 11371 28273
rect 11427 28243 11443 28273
rect 11495 28243 11515 28273
rect 11563 28243 11587 28273
rect 11631 28243 11659 28273
rect 11699 28243 11731 28273
rect 11223 28239 11257 28243
rect 11291 28239 11325 28243
rect 11359 28239 11393 28243
rect 11427 28239 11461 28243
rect 11495 28239 11529 28243
rect 11563 28239 11597 28243
rect 11631 28239 11665 28243
rect 11699 28239 11733 28243
rect 11767 28239 11801 28273
rect 11837 28243 11869 28273
rect 11909 28243 11937 28273
rect 11981 28243 12005 28273
rect 12053 28243 12073 28273
rect 12125 28243 12141 28273
rect 12197 28243 12209 28273
rect 12269 28243 12277 28273
rect 12341 28243 12345 28273
rect 11835 28239 11869 28243
rect 11903 28239 11937 28243
rect 11971 28239 12005 28243
rect 12039 28239 12073 28243
rect 12107 28239 12141 28243
rect 12175 28239 12209 28243
rect 12243 28239 12277 28243
rect 12311 28239 12345 28243
rect 12413 28273 12451 28277
rect 12485 28273 12523 28277
rect 12379 28239 12413 28243
rect 12447 28243 12451 28273
rect 12515 28243 12523 28273
rect 12557 28243 12832 28277
rect 12447 28239 12481 28243
rect 12515 28239 12832 28243
rect 2148 28203 12832 28239
rect 2148 28169 2479 28203
rect 2519 28169 2551 28203
rect 2587 28169 2621 28203
rect 2657 28169 2689 28203
rect 2729 28169 2757 28203
rect 2801 28169 2825 28203
rect 2873 28169 2893 28203
rect 2945 28169 2961 28203
rect 3017 28169 3029 28203
rect 3089 28169 3097 28203
rect 3161 28169 3165 28203
rect 3267 28169 3271 28203
rect 3335 28169 3343 28203
rect 3403 28169 3415 28203
rect 3471 28169 3487 28203
rect 3539 28169 3559 28203
rect 3607 28169 3631 28203
rect 3675 28169 3703 28203
rect 3743 28169 3775 28203
rect 3811 28169 3845 28203
rect 3881 28169 3913 28203
rect 3953 28169 3981 28203
rect 4025 28169 4049 28203
rect 4097 28169 4117 28203
rect 4169 28169 4185 28203
rect 4241 28169 4253 28203
rect 4313 28169 4321 28203
rect 4385 28169 4389 28203
rect 4491 28169 4495 28203
rect 4559 28169 4567 28203
rect 4627 28169 4639 28203
rect 4695 28169 4711 28203
rect 4763 28169 4783 28203
rect 4831 28169 4855 28203
rect 4899 28169 4927 28203
rect 4967 28169 4999 28203
rect 5035 28169 5069 28203
rect 5105 28169 5137 28203
rect 5177 28169 5205 28203
rect 5249 28169 5273 28203
rect 5321 28169 5341 28203
rect 5393 28169 5409 28203
rect 5465 28169 5477 28203
rect 5537 28169 5545 28203
rect 5609 28169 5613 28203
rect 5715 28169 5719 28203
rect 5783 28169 5791 28203
rect 5851 28169 5863 28203
rect 5919 28169 5935 28203
rect 5987 28169 6007 28203
rect 6055 28169 6079 28203
rect 6123 28169 6151 28203
rect 6191 28169 6223 28203
rect 6259 28169 6293 28203
rect 6329 28169 6361 28203
rect 6401 28169 6429 28203
rect 6473 28169 6497 28203
rect 6545 28169 6565 28203
rect 6617 28169 6633 28203
rect 6689 28169 6701 28203
rect 6761 28169 6769 28203
rect 6833 28169 6837 28203
rect 6939 28169 6943 28203
rect 7007 28169 7015 28203
rect 7075 28169 7087 28203
rect 7143 28169 7159 28203
rect 7211 28169 7231 28203
rect 7279 28169 7303 28203
rect 7347 28169 7375 28203
rect 7415 28169 7447 28203
rect 7483 28169 7517 28203
rect 7553 28169 7585 28203
rect 7625 28169 7653 28203
rect 7697 28169 7721 28203
rect 7769 28169 7789 28203
rect 7841 28169 7857 28203
rect 7913 28169 7925 28203
rect 7985 28169 7993 28203
rect 8057 28169 8061 28203
rect 8163 28169 8167 28203
rect 8231 28169 8239 28203
rect 8299 28169 8311 28203
rect 8367 28169 8383 28203
rect 8435 28169 8455 28203
rect 8503 28169 8527 28203
rect 8571 28169 8599 28203
rect 8639 28169 8671 28203
rect 8707 28169 8741 28203
rect 8777 28169 8809 28203
rect 8849 28169 8877 28203
rect 8921 28169 8945 28203
rect 8993 28169 9013 28203
rect 9065 28169 9081 28203
rect 9137 28169 9149 28203
rect 9209 28169 9217 28203
rect 9281 28169 9285 28203
rect 9387 28169 9391 28203
rect 9455 28169 9463 28203
rect 9523 28169 9535 28203
rect 9591 28169 9607 28203
rect 9659 28169 9679 28203
rect 9727 28169 9751 28203
rect 9795 28169 9823 28203
rect 9863 28169 9895 28203
rect 9931 28169 9965 28203
rect 10001 28169 10033 28203
rect 10073 28169 10101 28203
rect 10145 28169 10169 28203
rect 10217 28169 10237 28203
rect 10289 28169 10305 28203
rect 10361 28169 10373 28203
rect 10433 28169 10441 28203
rect 10505 28169 10509 28203
rect 10611 28169 10615 28203
rect 10679 28169 10687 28203
rect 10747 28169 10759 28203
rect 10815 28169 10831 28203
rect 10883 28169 10903 28203
rect 10951 28169 10975 28203
rect 11019 28169 11047 28203
rect 11087 28169 11119 28203
rect 11155 28169 11189 28203
rect 11225 28169 11257 28203
rect 11297 28169 11325 28203
rect 11369 28169 11393 28203
rect 11441 28169 11461 28203
rect 11513 28169 11529 28203
rect 11585 28169 11597 28203
rect 11657 28169 11665 28203
rect 11729 28169 11733 28203
rect 11835 28169 11839 28203
rect 11903 28169 11911 28203
rect 11971 28169 11983 28203
rect 12039 28169 12055 28203
rect 12107 28169 12127 28203
rect 12175 28169 12199 28203
rect 12243 28169 12271 28203
rect 12311 28169 12343 28203
rect 12379 28169 12413 28203
rect 12449 28169 12481 28203
rect 12521 28169 12832 28203
rect 2148 28104 2410 28169
rect 2148 28064 2376 28104
rect 12590 28104 12832 28169
rect 2148 28032 2410 28064
rect 2148 27996 2376 28032
rect 2148 27962 2410 27996
rect 2148 27926 2376 27962
rect 2148 27894 2410 27926
rect 2148 27854 2376 27894
rect 2496 28064 12504 28067
rect 2496 28032 2519 28064
rect 12481 28032 12504 28064
rect 2496 27926 2515 28032
rect 12485 27926 12504 28032
rect 2496 27894 2519 27926
rect 12481 27894 12504 27926
rect 2496 27891 12504 27894
rect 12624 28064 12832 28104
rect 12590 28032 12832 28064
rect 12624 27996 12832 28032
rect 12590 27962 12832 27996
rect 12624 27926 12832 27962
rect 12590 27894 12832 27926
rect 2148 27789 2410 27854
rect 12624 27854 12832 27894
rect 12590 27789 12832 27854
rect 2148 27717 2479 27789
rect 2148 27683 2443 27717
rect 2477 27683 2479 27717
rect 12521 27717 12832 27789
rect 12521 27683 12523 27717
rect 12557 27683 12832 27717
rect 2148 27569 12832 27683
rect 1651 27460 1718 27517
rect 1968 27464 2085 27517
rect 12915 27517 12945 28435
rect 13319 27517 13349 28435
rect 12915 27464 13023 27517
rect 1968 27460 13023 27464
rect 1651 27453 13023 27460
rect 13273 27453 13349 27517
rect 1651 27434 13349 27453
rect 1651 27347 2111 27434
rect 12889 27347 13349 27434
rect 1651 27097 1977 27347
rect 13027 27097 13349 27347
rect 1651 27060 2111 27097
rect 12889 27060 13349 27097
rect 1651 27030 13349 27060
rect 13761 28909 13801 28962
rect 13835 28909 13879 28962
rect 13761 28894 13879 28909
rect 13761 28837 13801 28894
rect 13835 28837 13879 28894
rect 13761 28826 13879 28837
rect 13761 28765 13801 28826
rect 13835 28765 13879 28826
rect 13761 28758 13879 28765
rect 13761 28724 13801 28758
rect 13835 28724 13879 28758
rect 13761 28690 13879 28724
rect 13761 28656 13801 28690
rect 13835 28656 13879 28690
rect 13761 28622 13879 28656
rect 13761 28588 13801 28622
rect 13835 28588 13879 28622
rect 13761 28554 13879 28588
rect 13761 28520 13801 28554
rect 13835 28520 13879 28554
rect 13761 28486 13879 28520
rect 13761 28452 13801 28486
rect 13835 28452 13879 28486
rect 13761 28418 13879 28452
rect 13761 28384 13801 28418
rect 13835 28384 13879 28418
rect 13761 28350 13879 28384
rect 13761 28316 13801 28350
rect 13835 28316 13879 28350
rect 13761 28282 13879 28316
rect 13761 28248 13801 28282
rect 13835 28248 13879 28282
rect 13761 28214 13879 28248
rect 13761 28180 13801 28214
rect 13835 28180 13879 28214
rect 13761 28146 13879 28180
rect 13761 28112 13801 28146
rect 13835 28112 13879 28146
rect 13761 28078 13879 28112
rect 13761 28044 13801 28078
rect 13835 28044 13879 28078
rect 13761 28010 13879 28044
rect 13761 27976 13801 28010
rect 13835 27976 13879 28010
rect 13761 27942 13879 27976
rect 13761 27908 13801 27942
rect 13835 27908 13879 27942
rect 13761 27874 13879 27908
rect 13761 27840 13801 27874
rect 13835 27840 13879 27874
rect 13761 27806 13879 27840
rect 13761 27772 13801 27806
rect 13835 27772 13879 27806
rect 13761 27738 13879 27772
rect 13761 27704 13801 27738
rect 13835 27704 13879 27738
rect 13761 27670 13879 27704
rect 13761 27636 13801 27670
rect 13835 27636 13879 27670
rect 13761 27602 13879 27636
rect 13761 27568 13801 27602
rect 13835 27568 13879 27602
rect 13761 27534 13879 27568
rect 13761 27500 13801 27534
rect 13835 27500 13879 27534
rect 13761 27466 13879 27500
rect 13761 27432 13801 27466
rect 13835 27432 13879 27466
rect 13761 27398 13879 27432
rect 13761 27364 13801 27398
rect 13835 27364 13879 27398
rect 13761 27330 13879 27364
rect 13761 27296 13801 27330
rect 13835 27296 13879 27330
rect 13761 27262 13879 27296
rect 13761 27228 13801 27262
rect 13835 27228 13879 27262
rect 13761 27194 13879 27228
rect 13761 27160 13801 27194
rect 13835 27160 13879 27194
rect 13761 27126 13879 27160
rect 13761 27092 13801 27126
rect 13835 27092 13879 27126
rect 13761 27058 13879 27092
rect 1111 27007 1229 27029
rect 1111 26961 1153 27007
rect 1187 26961 1229 27007
rect 1111 26935 1229 26961
rect 1111 26893 1153 26935
rect 1187 26893 1229 26935
rect 1111 26863 1229 26893
rect 1111 26825 1153 26863
rect 1187 26825 1229 26863
rect 1111 26791 1229 26825
rect 1111 26757 1153 26791
rect 1187 26757 1229 26791
rect 1111 26723 1229 26757
rect 1111 26685 1153 26723
rect 1187 26685 1229 26723
rect 1111 26655 1229 26685
rect 1111 26613 1153 26655
rect 1187 26613 1229 26655
rect 13761 27024 13801 27058
rect 13835 27024 13879 27058
rect 13761 26990 13879 27024
rect 13761 26956 13801 26990
rect 13835 26956 13879 26990
rect 13761 26922 13879 26956
rect 13761 26888 13801 26922
rect 13835 26888 13879 26922
rect 13761 26854 13879 26888
rect 13761 26820 13801 26854
rect 13835 26820 13879 26854
rect 13761 26786 13879 26820
rect 13761 26752 13801 26786
rect 13835 26752 13879 26786
rect 13761 26718 13879 26752
rect 13761 26684 13801 26718
rect 13835 26684 13879 26718
rect 13761 26650 13879 26684
rect 13761 26626 13801 26650
rect 1111 26587 1229 26613
rect 1111 26541 1153 26587
rect 1187 26541 1229 26587
rect 1111 26519 1229 26541
rect 1111 26469 1153 26519
rect 1187 26469 1229 26519
rect 1111 26451 1229 26469
rect 1111 26397 1153 26451
rect 1187 26397 1229 26451
rect 1111 26383 1229 26397
rect 1111 26325 1153 26383
rect 1187 26325 1229 26383
rect 1111 26315 1229 26325
rect 1111 26253 1153 26315
rect 1187 26253 1229 26315
rect 1111 26247 1229 26253
rect 1111 26181 1153 26247
rect 1187 26181 1229 26247
rect 1111 26179 1229 26181
rect 1111 26145 1153 26179
rect 1187 26145 1229 26179
rect 1111 26143 1229 26145
rect 1111 26077 1153 26143
rect 1187 26077 1229 26143
rect 1111 26071 1229 26077
rect 1111 26009 1153 26071
rect 1187 26009 1229 26071
rect 1111 25999 1229 26009
rect 1111 25941 1153 25999
rect 1187 25941 1229 25999
rect 1111 25927 1229 25941
rect 1111 25873 1153 25927
rect 1187 25873 1229 25927
rect 1111 25855 1229 25873
rect 1111 25805 1153 25855
rect 1187 25805 1229 25855
rect 1111 25783 1229 25805
rect 1111 25737 1153 25783
rect 1187 25737 1229 25783
rect 1111 25711 1229 25737
rect 1111 25669 1153 25711
rect 1187 25669 1229 25711
rect 1111 25639 1229 25669
rect 1111 25601 1153 25639
rect 1187 25601 1229 25639
rect 1111 25567 1229 25601
rect 1111 25533 1153 25567
rect 1187 25533 1229 25567
rect 1111 25499 1229 25533
rect 1111 25461 1153 25499
rect 1187 25461 1229 25499
rect 1111 25431 1229 25461
rect 1111 25389 1153 25431
rect 1187 25389 1229 25431
rect 1111 25363 1229 25389
rect 1111 25317 1153 25363
rect 1187 25317 1229 25363
rect 1111 25295 1229 25317
rect 1111 25245 1153 25295
rect 1187 25245 1229 25295
rect 1111 25227 1229 25245
rect 1111 25173 1153 25227
rect 1187 25173 1229 25227
rect 1111 25159 1229 25173
rect 1111 25101 1153 25159
rect 1187 25101 1229 25159
rect 1111 25091 1229 25101
rect 1111 25029 1153 25091
rect 1187 25029 1229 25091
rect 1111 25023 1229 25029
rect 1111 24957 1153 25023
rect 1187 24957 1229 25023
rect 1111 24955 1229 24957
rect 1111 24921 1153 24955
rect 1187 24921 1229 24955
rect 1111 24919 1229 24921
rect 1111 24853 1153 24919
rect 1187 24853 1229 24919
rect 1111 24847 1229 24853
rect 1111 24785 1153 24847
rect 1187 24785 1229 24847
rect 1690 26616 13801 26626
rect 13835 26616 13879 26650
rect 1690 26585 13879 26616
rect 1690 26191 2251 26585
rect 12725 26582 13879 26585
rect 12725 26548 13801 26582
rect 13835 26548 13879 26582
rect 12725 26514 13879 26548
rect 12725 26480 13801 26514
rect 13835 26480 13879 26514
rect 12725 26446 13879 26480
rect 12725 26412 13801 26446
rect 13835 26412 13879 26446
rect 12725 26378 13879 26412
rect 12725 26344 13801 26378
rect 13835 26344 13879 26378
rect 12725 26310 13879 26344
rect 12725 26276 13801 26310
rect 13835 26276 13879 26310
rect 12725 26242 13879 26276
rect 12725 26208 13801 26242
rect 13835 26208 13879 26242
rect 12725 26191 13879 26208
rect 1690 26174 13879 26191
rect 1690 26140 13801 26174
rect 13835 26140 13879 26174
rect 1690 26106 13879 26140
rect 1690 26093 13801 26106
rect 1690 26087 2262 26093
rect 1690 25333 1748 26087
rect 2142 25333 2262 26087
rect 12704 26087 13801 26093
rect 2320 25909 12656 25979
rect 2320 25875 2473 25909
rect 2537 25875 2541 25909
rect 2643 25875 2647 25909
rect 2711 25875 2719 25909
rect 2779 25875 2791 25909
rect 2847 25875 2863 25909
rect 2915 25875 2935 25909
rect 2983 25875 3007 25909
rect 3051 25875 3079 25909
rect 3119 25875 3151 25909
rect 3187 25875 3221 25909
rect 3257 25875 3289 25909
rect 3329 25875 3357 25909
rect 3401 25875 3425 25909
rect 3473 25875 3493 25909
rect 3545 25875 3561 25909
rect 3617 25875 3629 25909
rect 3689 25875 3697 25909
rect 3761 25875 3765 25909
rect 3867 25875 3871 25909
rect 3935 25875 3943 25909
rect 4003 25875 4015 25909
rect 4071 25875 4087 25909
rect 4139 25875 4159 25909
rect 4207 25875 4231 25909
rect 4275 25875 4303 25909
rect 4343 25875 4375 25909
rect 4411 25875 4445 25909
rect 4481 25875 4513 25909
rect 4553 25875 4581 25909
rect 4625 25875 4649 25909
rect 4697 25875 4717 25909
rect 4769 25875 4785 25909
rect 4841 25875 4853 25909
rect 4913 25875 4921 25909
rect 4985 25875 4989 25909
rect 5091 25875 5095 25909
rect 5159 25875 5167 25909
rect 5227 25875 5239 25909
rect 5295 25875 5311 25909
rect 5363 25875 5383 25909
rect 5431 25875 5455 25909
rect 5499 25875 5527 25909
rect 5567 25875 5599 25909
rect 5635 25875 5669 25909
rect 5705 25875 5737 25909
rect 5777 25875 5805 25909
rect 5849 25875 5873 25909
rect 5921 25875 5941 25909
rect 5993 25875 6009 25909
rect 6065 25875 6077 25909
rect 6137 25875 6145 25909
rect 6209 25875 6213 25909
rect 6315 25875 6319 25909
rect 6383 25875 6391 25909
rect 6451 25875 6463 25909
rect 6519 25875 6535 25909
rect 6587 25875 6607 25909
rect 6655 25875 6679 25909
rect 6723 25875 6751 25909
rect 6791 25875 6823 25909
rect 6859 25875 6893 25909
rect 6929 25875 6961 25909
rect 7001 25875 7029 25909
rect 7073 25875 7097 25909
rect 7145 25875 7165 25909
rect 7217 25875 7233 25909
rect 7289 25875 7301 25909
rect 7361 25875 7369 25909
rect 7433 25875 7437 25909
rect 7539 25875 7543 25909
rect 7607 25875 7615 25909
rect 7675 25875 7687 25909
rect 7743 25875 7759 25909
rect 7811 25875 7831 25909
rect 7879 25875 7903 25909
rect 7947 25875 7975 25909
rect 8015 25875 8047 25909
rect 8083 25875 8117 25909
rect 8153 25875 8185 25909
rect 8225 25875 8253 25909
rect 8297 25875 8321 25909
rect 8369 25875 8389 25909
rect 8441 25875 8457 25909
rect 8513 25875 8525 25909
rect 8585 25875 8593 25909
rect 8657 25875 8661 25909
rect 8763 25875 8767 25909
rect 8831 25875 8839 25909
rect 8899 25875 8911 25909
rect 8967 25875 8983 25909
rect 9035 25875 9055 25909
rect 9103 25875 9127 25909
rect 9171 25875 9199 25909
rect 9239 25875 9271 25909
rect 9307 25875 9341 25909
rect 9377 25875 9409 25909
rect 9449 25875 9477 25909
rect 9521 25875 9545 25909
rect 9593 25875 9613 25909
rect 9665 25875 9681 25909
rect 9737 25875 9749 25909
rect 9809 25875 9817 25909
rect 9881 25875 9885 25909
rect 9987 25875 9991 25909
rect 10055 25875 10063 25909
rect 10123 25875 10135 25909
rect 10191 25875 10207 25909
rect 10259 25875 10279 25909
rect 10327 25875 10351 25909
rect 10395 25875 10423 25909
rect 10463 25875 10495 25909
rect 10531 25875 10565 25909
rect 10601 25875 10633 25909
rect 10673 25875 10701 25909
rect 10745 25875 10769 25909
rect 10817 25875 10837 25909
rect 10889 25875 10905 25909
rect 10961 25875 10973 25909
rect 11033 25875 11041 25909
rect 11105 25875 11109 25909
rect 11211 25875 11215 25909
rect 11279 25875 11287 25909
rect 11347 25875 11359 25909
rect 11415 25875 11431 25909
rect 11483 25875 11503 25909
rect 11551 25875 11575 25909
rect 11619 25875 11647 25909
rect 11687 25875 11719 25909
rect 11755 25875 11789 25909
rect 11825 25875 11857 25909
rect 11897 25875 11925 25909
rect 11969 25875 11993 25909
rect 12041 25875 12061 25909
rect 12113 25875 12129 25909
rect 12185 25875 12197 25909
rect 12257 25875 12265 25909
rect 12329 25875 12333 25909
rect 12435 25875 12439 25909
rect 12503 25875 12656 25909
rect 2320 25826 2420 25875
rect 2320 25762 2386 25826
rect 12556 25826 12656 25875
rect 2320 25758 2420 25762
rect 2320 25656 2386 25758
rect 2320 25652 2420 25656
rect 2320 25588 2386 25652
rect 2484 25792 12492 25795
rect 2484 25760 2507 25792
rect 12469 25760 12492 25792
rect 2484 25654 2503 25760
rect 12473 25654 12492 25760
rect 2484 25622 2507 25654
rect 12469 25622 12492 25654
rect 2484 25619 12492 25622
rect 12590 25762 12656 25826
rect 12556 25758 12656 25762
rect 12590 25656 12656 25758
rect 12556 25652 12656 25656
rect 2320 25539 2420 25588
rect 12590 25588 12656 25652
rect 12556 25539 12656 25588
rect 2320 25505 2473 25539
rect 2537 25505 2541 25539
rect 2643 25505 2647 25539
rect 2711 25505 2719 25539
rect 2779 25505 2791 25539
rect 2847 25505 2863 25539
rect 2915 25505 2935 25539
rect 2983 25505 3007 25539
rect 3051 25505 3079 25539
rect 3119 25505 3151 25539
rect 3187 25505 3221 25539
rect 3257 25505 3289 25539
rect 3329 25505 3357 25539
rect 3401 25505 3425 25539
rect 3473 25505 3493 25539
rect 3545 25505 3561 25539
rect 3617 25505 3629 25539
rect 3689 25505 3697 25539
rect 3761 25505 3765 25539
rect 3867 25505 3871 25539
rect 3935 25505 3943 25539
rect 4003 25505 4015 25539
rect 4071 25505 4087 25539
rect 4139 25505 4159 25539
rect 4207 25505 4231 25539
rect 4275 25505 4303 25539
rect 4343 25505 4375 25539
rect 4411 25505 4445 25539
rect 4481 25505 4513 25539
rect 4553 25505 4581 25539
rect 4625 25505 4649 25539
rect 4697 25505 4717 25539
rect 4769 25505 4785 25539
rect 4841 25505 4853 25539
rect 4913 25505 4921 25539
rect 4985 25505 4989 25539
rect 5091 25505 5095 25539
rect 5159 25505 5167 25539
rect 5227 25505 5239 25539
rect 5295 25505 5311 25539
rect 5363 25505 5383 25539
rect 5431 25505 5455 25539
rect 5499 25505 5527 25539
rect 5567 25505 5599 25539
rect 5635 25505 5669 25539
rect 5705 25505 5737 25539
rect 5777 25505 5805 25539
rect 5849 25505 5873 25539
rect 5921 25505 5941 25539
rect 5993 25505 6009 25539
rect 6065 25505 6077 25539
rect 6137 25505 6145 25539
rect 6209 25505 6213 25539
rect 6315 25505 6319 25539
rect 6383 25505 6391 25539
rect 6451 25505 6463 25539
rect 6519 25505 6535 25539
rect 6587 25505 6607 25539
rect 6655 25505 6679 25539
rect 6723 25505 6751 25539
rect 6791 25505 6823 25539
rect 6859 25505 6893 25539
rect 6929 25505 6961 25539
rect 7001 25505 7029 25539
rect 7073 25505 7097 25539
rect 7145 25505 7165 25539
rect 7217 25505 7233 25539
rect 7289 25505 7301 25539
rect 7361 25505 7369 25539
rect 7433 25505 7437 25539
rect 7539 25505 7543 25539
rect 7607 25505 7615 25539
rect 7675 25505 7687 25539
rect 7743 25505 7759 25539
rect 7811 25505 7831 25539
rect 7879 25505 7903 25539
rect 7947 25505 7975 25539
rect 8015 25505 8047 25539
rect 8083 25505 8117 25539
rect 8153 25505 8185 25539
rect 8225 25505 8253 25539
rect 8297 25505 8321 25539
rect 8369 25505 8389 25539
rect 8441 25505 8457 25539
rect 8513 25505 8525 25539
rect 8585 25505 8593 25539
rect 8657 25505 8661 25539
rect 8763 25505 8767 25539
rect 8831 25505 8839 25539
rect 8899 25505 8911 25539
rect 8967 25505 8983 25539
rect 9035 25505 9055 25539
rect 9103 25505 9127 25539
rect 9171 25505 9199 25539
rect 9239 25505 9271 25539
rect 9307 25505 9341 25539
rect 9377 25505 9409 25539
rect 9449 25505 9477 25539
rect 9521 25505 9545 25539
rect 9593 25505 9613 25539
rect 9665 25505 9681 25539
rect 9737 25505 9749 25539
rect 9809 25505 9817 25539
rect 9881 25505 9885 25539
rect 9987 25505 9991 25539
rect 10055 25505 10063 25539
rect 10123 25505 10135 25539
rect 10191 25505 10207 25539
rect 10259 25505 10279 25539
rect 10327 25505 10351 25539
rect 10395 25505 10423 25539
rect 10463 25505 10495 25539
rect 10531 25505 10565 25539
rect 10601 25505 10633 25539
rect 10673 25505 10701 25539
rect 10745 25505 10769 25539
rect 10817 25505 10837 25539
rect 10889 25505 10905 25539
rect 10961 25505 10973 25539
rect 11033 25505 11041 25539
rect 11105 25505 11109 25539
rect 11211 25505 11215 25539
rect 11279 25505 11287 25539
rect 11347 25505 11359 25539
rect 11415 25505 11431 25539
rect 11483 25505 11503 25539
rect 11551 25505 11575 25539
rect 11619 25505 11647 25539
rect 11687 25505 11719 25539
rect 11755 25505 11789 25539
rect 11825 25505 11857 25539
rect 11897 25505 11925 25539
rect 11969 25505 11993 25539
rect 12041 25505 12061 25539
rect 12113 25505 12129 25539
rect 12185 25505 12197 25539
rect 12257 25505 12265 25539
rect 12329 25505 12333 25539
rect 12435 25505 12439 25539
rect 12503 25505 12656 25539
rect 2320 25441 12656 25505
rect 1690 25326 2262 25333
rect 12704 25333 12834 26087
rect 13228 26072 13801 26087
rect 13835 26072 13879 26106
rect 13228 26038 13879 26072
rect 13228 26004 13801 26038
rect 13835 26004 13879 26038
rect 13228 25970 13879 26004
rect 13228 25936 13801 25970
rect 13835 25936 13879 25970
rect 13228 25902 13879 25936
rect 13228 25868 13801 25902
rect 13835 25868 13879 25902
rect 13228 25834 13879 25868
rect 13228 25800 13801 25834
rect 13835 25800 13879 25834
rect 13228 25766 13879 25800
rect 13228 25732 13801 25766
rect 13835 25732 13879 25766
rect 13228 25698 13879 25732
rect 13228 25664 13801 25698
rect 13835 25664 13879 25698
rect 13228 25630 13879 25664
rect 13228 25596 13801 25630
rect 13835 25596 13879 25630
rect 13228 25562 13879 25596
rect 13228 25528 13801 25562
rect 13835 25528 13879 25562
rect 13228 25494 13879 25528
rect 13228 25460 13801 25494
rect 13835 25460 13879 25494
rect 13228 25426 13879 25460
rect 13228 25392 13801 25426
rect 13835 25392 13879 25426
rect 13228 25358 13879 25392
rect 13228 25333 13801 25358
rect 12704 25326 13801 25333
rect 1690 25324 13801 25326
rect 13835 25324 13879 25358
rect 1690 25290 13879 25324
rect 1690 25256 13801 25290
rect 13835 25256 13879 25290
rect 1690 25229 13879 25256
rect 1690 24835 2251 25229
rect 12725 25222 13879 25229
rect 12725 25188 13801 25222
rect 13835 25188 13879 25222
rect 12725 25154 13879 25188
rect 12725 25120 13801 25154
rect 13835 25120 13879 25154
rect 12725 25086 13879 25120
rect 12725 25052 13801 25086
rect 13835 25052 13879 25086
rect 12725 25018 13879 25052
rect 12725 24984 13801 25018
rect 13835 24984 13879 25018
rect 12725 24950 13879 24984
rect 12725 24916 13801 24950
rect 13835 24916 13879 24950
rect 12725 24882 13879 24916
rect 12725 24848 13801 24882
rect 13835 24848 13879 24882
rect 12725 24835 13879 24848
rect 1690 24814 13879 24835
rect 1690 24793 13801 24814
rect 1111 24775 1229 24785
rect 1111 24717 1153 24775
rect 1187 24717 1229 24775
rect 1111 24703 1229 24717
rect 1111 24649 1153 24703
rect 1187 24649 1229 24703
rect 1111 24631 1229 24649
rect 1111 24581 1153 24631
rect 1187 24581 1229 24631
rect 1111 24559 1229 24581
rect 1111 24513 1153 24559
rect 1187 24513 1229 24559
rect 1111 24487 1229 24513
rect 1111 24445 1153 24487
rect 1187 24445 1229 24487
rect 1111 24415 1229 24445
rect 1111 24377 1153 24415
rect 1187 24377 1229 24415
rect 1111 24343 1229 24377
rect 1111 24309 1153 24343
rect 1187 24309 1229 24343
rect 1111 24275 1229 24309
rect 1111 24237 1153 24275
rect 1187 24237 1229 24275
rect 1111 24207 1229 24237
rect 1111 24165 1153 24207
rect 1187 24165 1229 24207
rect 1111 24139 1229 24165
rect 1111 24093 1153 24139
rect 1187 24093 1229 24139
rect 1111 24071 1229 24093
rect 1111 24021 1153 24071
rect 1187 24021 1229 24071
rect 1111 24003 1229 24021
rect 1111 23949 1153 24003
rect 1187 23949 1229 24003
rect 1111 23935 1229 23949
rect 1111 23877 1153 23935
rect 1187 23877 1229 23935
rect 1111 23867 1229 23877
rect 1111 23805 1153 23867
rect 1187 23805 1229 23867
rect 1111 23799 1229 23805
rect 1111 23733 1153 23799
rect 1187 23733 1229 23799
rect 1111 23731 1229 23733
rect 1111 23697 1153 23731
rect 1187 23697 1229 23731
rect 1111 23695 1229 23697
rect 1111 23629 1153 23695
rect 1187 23629 1229 23695
rect 1111 23623 1229 23629
rect 1111 23561 1153 23623
rect 1187 23561 1229 23623
rect 1111 23551 1229 23561
rect 1111 23493 1153 23551
rect 1187 23493 1229 23551
rect 1111 23479 1229 23493
rect 1111 23425 1153 23479
rect 1187 23425 1229 23479
rect 1111 23407 1229 23425
rect 1111 23357 1153 23407
rect 1187 23357 1229 23407
rect 1111 23335 1229 23357
rect 1111 23289 1153 23335
rect 1187 23289 1229 23335
rect 1111 23263 1229 23289
rect 1111 23221 1153 23263
rect 1187 23221 1229 23263
rect 1111 23191 1229 23221
rect 1111 23153 1153 23191
rect 1187 23153 1229 23191
rect 1111 23119 1229 23153
rect 1111 23085 1153 23119
rect 1187 23085 1229 23119
rect 1111 23051 1229 23085
rect 1111 23013 1153 23051
rect 1187 23013 1229 23051
rect 1111 22983 1229 23013
rect 1111 22941 1153 22983
rect 1187 22941 1229 22983
rect 1111 22915 1229 22941
rect 1111 22869 1153 22915
rect 1187 22869 1229 22915
rect 1111 22847 1229 22869
rect 1111 22797 1153 22847
rect 1187 22797 1229 22847
rect 1111 22779 1229 22797
rect 1111 22725 1153 22779
rect 1187 22725 1229 22779
rect 1111 22711 1229 22725
rect 1111 22653 1153 22711
rect 1187 22653 1229 22711
rect 1111 22643 1229 22653
rect 1111 22581 1153 22643
rect 1187 22581 1229 22643
rect 1111 22575 1229 22581
rect 1111 22509 1153 22575
rect 1187 22509 1229 22575
rect 1111 22507 1229 22509
rect 1111 22473 1153 22507
rect 1187 22473 1229 22507
rect 1111 22471 1229 22473
rect 1111 22405 1153 22471
rect 1187 22405 1229 22471
rect 1111 22399 1229 22405
rect 1111 22337 1153 22399
rect 1187 22337 1229 22399
rect 1111 22327 1229 22337
rect 1111 22269 1153 22327
rect 1187 22269 1229 22327
rect 1111 22255 1229 22269
rect 1111 22201 1153 22255
rect 1187 22201 1229 22255
rect 1111 22183 1229 22201
rect 1111 22133 1153 22183
rect 1187 22133 1229 22183
rect 1111 22111 1229 22133
rect 1111 22065 1153 22111
rect 1187 22065 1229 22111
rect 1111 22039 1229 22065
rect 1111 21997 1153 22039
rect 1187 21997 1229 22039
rect 1111 21967 1229 21997
rect 1111 21929 1153 21967
rect 1187 21929 1229 21967
rect 1111 21895 1229 21929
rect 1111 21861 1153 21895
rect 1187 21861 1229 21895
rect 1111 21827 1229 21861
rect 1111 21789 1153 21827
rect 1187 21789 1229 21827
rect 1111 21759 1229 21789
rect 1111 21717 1153 21759
rect 1187 21717 1229 21759
rect 1111 21691 1229 21717
rect 1111 21645 1153 21691
rect 1187 21645 1229 21691
rect 1111 21623 1229 21645
rect 1111 21573 1153 21623
rect 1187 21573 1229 21623
rect 1111 21555 1229 21573
rect 1111 21501 1153 21555
rect 1187 21501 1229 21555
rect 1111 21487 1229 21501
rect 1111 21429 1153 21487
rect 1187 21429 1229 21487
rect 1111 21419 1229 21429
rect 1111 21357 1153 21419
rect 1187 21357 1229 21419
rect 1111 21351 1229 21357
rect 1111 21285 1153 21351
rect 1187 21285 1229 21351
rect 1111 21283 1229 21285
rect 1111 21249 1153 21283
rect 1187 21249 1229 21283
rect 1111 21247 1229 21249
rect 1111 21181 1153 21247
rect 1187 21181 1229 21247
rect 1111 21175 1229 21181
rect 1111 21113 1153 21175
rect 1187 21113 1229 21175
rect 1111 21103 1229 21113
rect 1111 21045 1153 21103
rect 1187 21045 1229 21103
rect 1111 21031 1229 21045
rect 1111 20977 1153 21031
rect 1187 20977 1229 21031
rect 1111 20959 1229 20977
rect 1111 20909 1153 20959
rect 1187 20909 1229 20959
rect 1111 20887 1229 20909
rect 1111 20841 1153 20887
rect 1187 20841 1229 20887
rect 1111 20815 1229 20841
rect 1111 20773 1153 20815
rect 1187 20773 1229 20815
rect 1111 20743 1229 20773
rect 1111 20705 1153 20743
rect 1187 20705 1229 20743
rect 1111 20671 1229 20705
rect 1111 20637 1153 20671
rect 1187 20637 1229 20671
rect 1111 20603 1229 20637
rect 1111 20565 1153 20603
rect 1187 20565 1229 20603
rect 1111 20535 1229 20565
rect 1111 20493 1153 20535
rect 1187 20493 1229 20535
rect 1111 20467 1229 20493
rect 1111 20421 1153 20467
rect 1187 20421 1229 20467
rect 1111 20399 1229 20421
rect 1111 20349 1153 20399
rect 1187 20349 1229 20399
rect 1111 20331 1229 20349
rect 1111 20277 1153 20331
rect 1187 20277 1229 20331
rect 1111 20263 1229 20277
rect 1111 20205 1153 20263
rect 1187 20205 1229 20263
rect 1111 20195 1229 20205
rect 1111 20133 1153 20195
rect 1187 20133 1229 20195
rect 1111 20127 1229 20133
rect 1111 20061 1153 20127
rect 1187 20061 1229 20127
rect 1111 20059 1229 20061
rect 1111 20025 1153 20059
rect 1187 20025 1229 20059
rect 1111 20023 1229 20025
rect 1111 19957 1153 20023
rect 1187 19957 1229 20023
rect 1111 19951 1229 19957
rect 1111 19889 1153 19951
rect 1187 19889 1229 19951
rect 1111 19879 1229 19889
rect 1111 19821 1153 19879
rect 1187 19821 1229 19879
rect 1111 19807 1229 19821
rect 1111 19753 1153 19807
rect 1187 19753 1229 19807
rect 1111 19735 1229 19753
rect 1111 19685 1153 19735
rect 1187 19685 1229 19735
rect 1111 19663 1229 19685
rect 1111 19617 1153 19663
rect 1187 19617 1229 19663
rect 1111 19591 1229 19617
rect 1111 19549 1153 19591
rect 1187 19549 1229 19591
rect 1111 19519 1229 19549
rect 1111 19481 1153 19519
rect 1187 19481 1229 19519
rect 1111 19447 1229 19481
rect 1111 19413 1153 19447
rect 1187 19413 1229 19447
rect 1111 19379 1229 19413
rect 1111 19341 1153 19379
rect 1187 19341 1229 19379
rect 1111 19311 1229 19341
rect 1111 19269 1153 19311
rect 1187 19269 1229 19311
rect 1111 19243 1229 19269
rect 1111 19197 1153 19243
rect 1187 19197 1229 19243
rect 1111 19175 1229 19197
rect 1111 19125 1153 19175
rect 1187 19125 1229 19175
rect 1111 19107 1229 19125
rect 1111 19053 1153 19107
rect 1187 19053 1229 19107
rect 1111 19039 1229 19053
rect 1111 18981 1153 19039
rect 1187 18981 1229 19039
rect 1111 18971 1229 18981
rect 1111 18909 1153 18971
rect 1187 18909 1229 18971
rect 1111 18903 1229 18909
rect 1111 18837 1153 18903
rect 1187 18837 1229 18903
rect 1111 18835 1229 18837
rect 1111 18801 1153 18835
rect 1187 18801 1229 18835
rect 1111 18799 1229 18801
rect 1111 18733 1153 18799
rect 1187 18733 1229 18799
rect 1111 18727 1229 18733
rect 1111 18665 1153 18727
rect 1187 18665 1229 18727
rect 1111 18655 1229 18665
rect 1111 18597 1153 18655
rect 1187 18597 1229 18655
rect 1111 18583 1229 18597
rect 1111 18529 1153 18583
rect 1187 18529 1229 18583
rect 1111 18511 1229 18529
rect 1111 18461 1153 18511
rect 1187 18461 1229 18511
rect 1111 18439 1229 18461
rect 1111 18393 1153 18439
rect 1187 18393 1229 18439
rect 1111 18367 1229 18393
rect 1111 18325 1153 18367
rect 1187 18325 1229 18367
rect 1111 18295 1229 18325
rect 1111 18257 1153 18295
rect 1187 18257 1229 18295
rect 1111 18223 1229 18257
rect 1111 18189 1153 18223
rect 1187 18189 1229 18223
rect 1111 18155 1229 18189
rect 1111 18117 1153 18155
rect 1187 18117 1229 18155
rect 1111 18087 1229 18117
rect 1111 18045 1153 18087
rect 1187 18045 1229 18087
rect 1111 18019 1229 18045
rect 1111 17973 1153 18019
rect 1187 17973 1229 18019
rect 1111 17951 1229 17973
rect 1111 17901 1153 17951
rect 1187 17901 1229 17951
rect 1111 17883 1229 17901
rect 1111 17829 1153 17883
rect 1187 17829 1229 17883
rect 1111 17815 1229 17829
rect 1111 17757 1153 17815
rect 1187 17757 1229 17815
rect 1111 17747 1229 17757
rect 1111 17685 1153 17747
rect 1187 17685 1229 17747
rect 1111 17679 1229 17685
rect 1111 17613 1153 17679
rect 1187 17613 1229 17679
rect 1111 17611 1229 17613
rect 1111 17577 1153 17611
rect 1187 17577 1229 17611
rect 1111 17575 1229 17577
rect 1111 17509 1153 17575
rect 1187 17509 1229 17575
rect 1111 17503 1229 17509
rect 1111 17441 1153 17503
rect 1187 17441 1229 17503
rect 1111 17431 1229 17441
rect 1111 17373 1153 17431
rect 1187 17373 1229 17431
rect 1111 17359 1229 17373
rect 1111 17305 1153 17359
rect 1187 17305 1229 17359
rect 1111 17287 1229 17305
rect 1111 17237 1153 17287
rect 1187 17237 1229 17287
rect 1111 17215 1229 17237
rect 1111 17169 1153 17215
rect 1187 17169 1229 17215
rect 1111 17143 1229 17169
rect 1111 17101 1153 17143
rect 1187 17101 1229 17143
rect 1111 17071 1229 17101
rect 1111 17033 1153 17071
rect 1187 17033 1229 17071
rect 1111 16999 1229 17033
rect 1111 16965 1153 16999
rect 1187 16965 1229 16999
rect 1111 16931 1229 16965
rect 1111 16893 1153 16931
rect 1187 16893 1229 16931
rect 1111 16863 1229 16893
rect 1111 16821 1153 16863
rect 1187 16821 1229 16863
rect 1111 16795 1229 16821
rect 1111 16749 1153 16795
rect 1187 16749 1229 16795
rect 1111 16727 1229 16749
rect 1111 16677 1153 16727
rect 1187 16677 1229 16727
rect 1111 16659 1229 16677
rect 1111 16605 1153 16659
rect 1187 16605 1229 16659
rect 1111 16591 1229 16605
rect 1111 16533 1153 16591
rect 1187 16533 1229 16591
rect 1111 16523 1229 16533
rect 1111 16461 1153 16523
rect 1187 16461 1229 16523
rect 1111 16455 1229 16461
rect 1111 16389 1153 16455
rect 1187 16389 1229 16455
rect 1111 16387 1229 16389
rect 1111 16353 1153 16387
rect 1187 16353 1229 16387
rect 1111 16351 1229 16353
rect 1111 16285 1153 16351
rect 1187 16285 1229 16351
rect 1111 16279 1229 16285
rect 1111 16217 1153 16279
rect 1187 16217 1229 16279
rect 1111 16207 1229 16217
rect 1111 16149 1153 16207
rect 1187 16149 1229 16207
rect 1111 16135 1229 16149
rect 1111 16081 1153 16135
rect 1187 16081 1229 16135
rect 1111 16063 1229 16081
rect 1111 16013 1153 16063
rect 1187 16013 1229 16063
rect 1111 15991 1229 16013
rect 1111 15945 1153 15991
rect 1187 15945 1229 15991
rect 1111 15919 1229 15945
rect 1111 15877 1153 15919
rect 1187 15877 1229 15919
rect 1111 15847 1229 15877
rect 1111 15809 1153 15847
rect 1187 15809 1229 15847
rect 1111 15775 1229 15809
rect 1111 15741 1153 15775
rect 1187 15741 1229 15775
rect 1111 15707 1229 15741
rect 1111 15669 1153 15707
rect 1187 15669 1229 15707
rect 1111 15639 1229 15669
rect 1111 15597 1153 15639
rect 1187 15597 1229 15639
rect 1111 15571 1229 15597
rect 1111 15525 1153 15571
rect 1187 15525 1229 15571
rect 1111 15503 1229 15525
rect 1111 15453 1153 15503
rect 1187 15453 1229 15503
rect 1111 15435 1229 15453
rect 1111 15381 1153 15435
rect 1187 15381 1229 15435
rect 1111 15332 1229 15381
rect 13761 24780 13801 24793
rect 13835 24780 13879 24814
rect 13761 24746 13879 24780
rect 13761 24712 13801 24746
rect 13835 24712 13879 24746
rect 13761 24678 13879 24712
rect 13761 24644 13801 24678
rect 13835 24644 13879 24678
rect 13761 24610 13879 24644
rect 13761 24576 13801 24610
rect 13835 24576 13879 24610
rect 13761 24542 13879 24576
rect 13761 24508 13801 24542
rect 13835 24508 13879 24542
rect 13761 24474 13879 24508
rect 13761 24440 13801 24474
rect 13835 24440 13879 24474
rect 13761 24406 13879 24440
rect 13761 24372 13801 24406
rect 13835 24372 13879 24406
rect 13761 24338 13879 24372
rect 13761 24304 13801 24338
rect 13835 24304 13879 24338
rect 13761 24270 13879 24304
rect 13761 24236 13801 24270
rect 13835 24236 13879 24270
rect 13761 24202 13879 24236
rect 13761 24168 13801 24202
rect 13835 24168 13879 24202
rect 13761 24134 13879 24168
rect 13761 24100 13801 24134
rect 13835 24100 13879 24134
rect 13761 24066 13879 24100
rect 13761 24032 13801 24066
rect 13835 24032 13879 24066
rect 13761 23998 13879 24032
rect 13761 23964 13801 23998
rect 13835 23964 13879 23998
rect 13761 23930 13879 23964
rect 13761 23896 13801 23930
rect 13835 23896 13879 23930
rect 13761 23862 13879 23896
rect 13761 23828 13801 23862
rect 13835 23828 13879 23862
rect 13761 23794 13879 23828
rect 13761 23760 13801 23794
rect 13835 23760 13879 23794
rect 13761 23726 13879 23760
rect 13761 23692 13801 23726
rect 13835 23692 13879 23726
rect 13761 23658 13879 23692
rect 13761 23624 13801 23658
rect 13835 23624 13879 23658
rect 13761 23590 13879 23624
rect 13761 23556 13801 23590
rect 13835 23556 13879 23590
rect 13761 23522 13879 23556
rect 13761 23488 13801 23522
rect 13835 23488 13879 23522
rect 13761 23454 13879 23488
rect 13761 23420 13801 23454
rect 13835 23420 13879 23454
rect 13761 23410 13879 23420
rect 13761 23352 13801 23410
rect 13835 23352 13879 23410
rect 13761 23338 13879 23352
rect 13761 23284 13801 23338
rect 13835 23284 13879 23338
rect 13761 23266 13879 23284
rect 13761 23216 13801 23266
rect 13835 23216 13879 23266
rect 13761 23194 13879 23216
rect 13761 23148 13801 23194
rect 13835 23148 13879 23194
rect 13761 23122 13879 23148
rect 13761 23080 13801 23122
rect 13835 23080 13879 23122
rect 13761 23050 13879 23080
rect 13761 23012 13801 23050
rect 13835 23012 13879 23050
rect 13761 22978 13879 23012
rect 13761 22944 13801 22978
rect 13835 22944 13879 22978
rect 13761 22910 13879 22944
rect 13761 22872 13801 22910
rect 13835 22872 13879 22910
rect 13761 22842 13879 22872
rect 13761 22800 13801 22842
rect 13835 22800 13879 22842
rect 13761 22774 13879 22800
rect 13761 22728 13801 22774
rect 13835 22728 13879 22774
rect 13761 22706 13879 22728
rect 13761 22656 13801 22706
rect 13835 22656 13879 22706
rect 13761 22638 13879 22656
rect 13761 22584 13801 22638
rect 13835 22584 13879 22638
rect 13761 22570 13879 22584
rect 13761 22512 13801 22570
rect 13835 22512 13879 22570
rect 13761 22502 13879 22512
rect 13761 22440 13801 22502
rect 13835 22440 13879 22502
rect 13761 22434 13879 22440
rect 13761 22368 13801 22434
rect 13835 22368 13879 22434
rect 13761 22366 13879 22368
rect 13761 22332 13801 22366
rect 13835 22332 13879 22366
rect 13761 22330 13879 22332
rect 13761 22264 13801 22330
rect 13835 22264 13879 22330
rect 13761 22258 13879 22264
rect 13761 22196 13801 22258
rect 13835 22196 13879 22258
rect 13761 22186 13879 22196
rect 13761 22128 13801 22186
rect 13835 22128 13879 22186
rect 13761 22114 13879 22128
rect 13761 22060 13801 22114
rect 13835 22060 13879 22114
rect 13761 22042 13879 22060
rect 13761 21992 13801 22042
rect 13835 21992 13879 22042
rect 13761 21970 13879 21992
rect 13761 21924 13801 21970
rect 13835 21924 13879 21970
rect 13761 21898 13879 21924
rect 13761 21856 13801 21898
rect 13835 21856 13879 21898
rect 13761 21826 13879 21856
rect 13761 21788 13801 21826
rect 13835 21788 13879 21826
rect 13761 21754 13879 21788
rect 13761 21720 13801 21754
rect 13835 21720 13879 21754
rect 13761 21686 13879 21720
rect 13761 21648 13801 21686
rect 13835 21648 13879 21686
rect 13761 21618 13879 21648
rect 13761 21576 13801 21618
rect 13835 21576 13879 21618
rect 13761 21550 13879 21576
rect 13761 21504 13801 21550
rect 13835 21504 13879 21550
rect 13761 21482 13879 21504
rect 13761 21432 13801 21482
rect 13835 21432 13879 21482
rect 13761 21414 13879 21432
rect 13761 21360 13801 21414
rect 13835 21360 13879 21414
rect 13761 21346 13879 21360
rect 13761 21288 13801 21346
rect 13835 21288 13879 21346
rect 13761 21278 13879 21288
rect 13761 21216 13801 21278
rect 13835 21216 13879 21278
rect 13761 21210 13879 21216
rect 13761 21144 13801 21210
rect 13835 21144 13879 21210
rect 13761 21142 13879 21144
rect 13761 21108 13801 21142
rect 13835 21108 13879 21142
rect 13761 21106 13879 21108
rect 13761 21040 13801 21106
rect 13835 21040 13879 21106
rect 13761 21034 13879 21040
rect 13761 20972 13801 21034
rect 13835 20972 13879 21034
rect 13761 20962 13879 20972
rect 13761 20904 13801 20962
rect 13835 20904 13879 20962
rect 13761 20890 13879 20904
rect 13761 20836 13801 20890
rect 13835 20836 13879 20890
rect 13761 20818 13879 20836
rect 13761 20768 13801 20818
rect 13835 20768 13879 20818
rect 13761 20746 13879 20768
rect 13761 20700 13801 20746
rect 13835 20700 13879 20746
rect 13761 20674 13879 20700
rect 13761 20632 13801 20674
rect 13835 20632 13879 20674
rect 13761 20602 13879 20632
rect 13761 20564 13801 20602
rect 13835 20564 13879 20602
rect 13761 20530 13879 20564
rect 13761 20496 13801 20530
rect 13835 20496 13879 20530
rect 13761 20462 13879 20496
rect 13761 20424 13801 20462
rect 13835 20424 13879 20462
rect 13761 20394 13879 20424
rect 13761 20352 13801 20394
rect 13835 20352 13879 20394
rect 13761 20326 13879 20352
rect 13761 20280 13801 20326
rect 13835 20280 13879 20326
rect 13761 20258 13879 20280
rect 13761 20208 13801 20258
rect 13835 20208 13879 20258
rect 13761 20190 13879 20208
rect 13761 20136 13801 20190
rect 13835 20136 13879 20190
rect 13761 20122 13879 20136
rect 13761 20064 13801 20122
rect 13835 20064 13879 20122
rect 13761 20054 13879 20064
rect 13761 19992 13801 20054
rect 13835 19992 13879 20054
rect 13761 19986 13879 19992
rect 13761 19920 13801 19986
rect 13835 19920 13879 19986
rect 13761 19918 13879 19920
rect 13761 19884 13801 19918
rect 13835 19884 13879 19918
rect 13761 19882 13879 19884
rect 13761 19816 13801 19882
rect 13835 19816 13879 19882
rect 13761 19810 13879 19816
rect 13761 19748 13801 19810
rect 13835 19748 13879 19810
rect 13761 19738 13879 19748
rect 13761 19680 13801 19738
rect 13835 19680 13879 19738
rect 13761 19666 13879 19680
rect 13761 19612 13801 19666
rect 13835 19612 13879 19666
rect 13761 19594 13879 19612
rect 13761 19544 13801 19594
rect 13835 19544 13879 19594
rect 13761 19522 13879 19544
rect 13761 19476 13801 19522
rect 13835 19476 13879 19522
rect 13761 19450 13879 19476
rect 13761 19408 13801 19450
rect 13835 19408 13879 19450
rect 13761 19378 13879 19408
rect 13761 19340 13801 19378
rect 13835 19340 13879 19378
rect 13761 19306 13879 19340
rect 13761 19272 13801 19306
rect 13835 19272 13879 19306
rect 13761 19238 13879 19272
rect 13761 19200 13801 19238
rect 13835 19200 13879 19238
rect 13761 19170 13879 19200
rect 13761 19128 13801 19170
rect 13835 19128 13879 19170
rect 13761 19102 13879 19128
rect 13761 19056 13801 19102
rect 13835 19056 13879 19102
rect 13761 19034 13879 19056
rect 13761 18984 13801 19034
rect 13835 18984 13879 19034
rect 13761 18966 13879 18984
rect 13761 18912 13801 18966
rect 13835 18912 13879 18966
rect 13761 18898 13879 18912
rect 13761 18840 13801 18898
rect 13835 18840 13879 18898
rect 13761 18830 13879 18840
rect 13761 18768 13801 18830
rect 13835 18768 13879 18830
rect 13761 18762 13879 18768
rect 13761 18696 13801 18762
rect 13835 18696 13879 18762
rect 13761 18694 13879 18696
rect 13761 18660 13801 18694
rect 13835 18660 13879 18694
rect 13761 18658 13879 18660
rect 13761 18592 13801 18658
rect 13835 18592 13879 18658
rect 13761 18586 13879 18592
rect 13761 18524 13801 18586
rect 13835 18524 13879 18586
rect 13761 18514 13879 18524
rect 13761 18456 13801 18514
rect 13835 18456 13879 18514
rect 13761 18442 13879 18456
rect 13761 18388 13801 18442
rect 13835 18388 13879 18442
rect 13761 18370 13879 18388
rect 13761 18320 13801 18370
rect 13835 18320 13879 18370
rect 13761 18298 13879 18320
rect 13761 18252 13801 18298
rect 13835 18252 13879 18298
rect 13761 18226 13879 18252
rect 13761 18184 13801 18226
rect 13835 18184 13879 18226
rect 13761 18154 13879 18184
rect 13761 18116 13801 18154
rect 13835 18116 13879 18154
rect 13761 18082 13879 18116
rect 13761 18048 13801 18082
rect 13835 18048 13879 18082
rect 13761 18014 13879 18048
rect 13761 17976 13801 18014
rect 13835 17976 13879 18014
rect 13761 17946 13879 17976
rect 13761 17904 13801 17946
rect 13835 17904 13879 17946
rect 13761 17878 13879 17904
rect 13761 17832 13801 17878
rect 13835 17832 13879 17878
rect 13761 17810 13879 17832
rect 13761 17760 13801 17810
rect 13835 17760 13879 17810
rect 13761 17742 13879 17760
rect 13761 17688 13801 17742
rect 13835 17688 13879 17742
rect 13761 17674 13879 17688
rect 13761 17616 13801 17674
rect 13835 17616 13879 17674
rect 13761 17606 13879 17616
rect 13761 17544 13801 17606
rect 13835 17544 13879 17606
rect 13761 17538 13879 17544
rect 13761 17472 13801 17538
rect 13835 17472 13879 17538
rect 13761 17470 13879 17472
rect 13761 17436 13801 17470
rect 13835 17436 13879 17470
rect 13761 17434 13879 17436
rect 13761 17368 13801 17434
rect 13835 17368 13879 17434
rect 13761 17362 13879 17368
rect 13761 17300 13801 17362
rect 13835 17300 13879 17362
rect 13761 17290 13879 17300
rect 13761 17232 13801 17290
rect 13835 17232 13879 17290
rect 13761 17218 13879 17232
rect 13761 17164 13801 17218
rect 13835 17164 13879 17218
rect 13761 17146 13879 17164
rect 13761 17096 13801 17146
rect 13835 17096 13879 17146
rect 13761 17074 13879 17096
rect 13761 17028 13801 17074
rect 13835 17028 13879 17074
rect 13761 17002 13879 17028
rect 13761 16960 13801 17002
rect 13835 16960 13879 17002
rect 13761 16930 13879 16960
rect 13761 16892 13801 16930
rect 13835 16892 13879 16930
rect 13761 16858 13879 16892
rect 13761 16824 13801 16858
rect 13835 16824 13879 16858
rect 13761 16790 13879 16824
rect 13761 16752 13801 16790
rect 13835 16752 13879 16790
rect 13761 16722 13879 16752
rect 13761 16680 13801 16722
rect 13835 16680 13879 16722
rect 13761 16654 13879 16680
rect 13761 16608 13801 16654
rect 13835 16608 13879 16654
rect 13761 16586 13879 16608
rect 13761 16536 13801 16586
rect 13835 16536 13879 16586
rect 13761 16518 13879 16536
rect 13761 16464 13801 16518
rect 13835 16464 13879 16518
rect 13761 16450 13879 16464
rect 13761 16392 13801 16450
rect 13835 16392 13879 16450
rect 13761 16382 13879 16392
rect 13761 16320 13801 16382
rect 13835 16320 13879 16382
rect 13761 16314 13879 16320
rect 13761 16248 13801 16314
rect 13835 16248 13879 16314
rect 13761 16246 13879 16248
rect 13761 16212 13801 16246
rect 13835 16212 13879 16246
rect 13761 16210 13879 16212
rect 13761 16144 13801 16210
rect 13835 16144 13879 16210
rect 13761 16138 13879 16144
rect 13761 16076 13801 16138
rect 13835 16076 13879 16138
rect 13761 16066 13879 16076
rect 13761 16008 13801 16066
rect 13835 16008 13879 16066
rect 13761 15994 13879 16008
rect 13761 15940 13801 15994
rect 13835 15940 13879 15994
rect 13761 15922 13879 15940
rect 13761 15872 13801 15922
rect 13835 15872 13879 15922
rect 13761 15850 13879 15872
rect 13761 15804 13801 15850
rect 13835 15804 13879 15850
rect 13761 15778 13879 15804
rect 13761 15736 13801 15778
rect 13835 15736 13879 15778
rect 13761 15706 13879 15736
rect 13761 15668 13801 15706
rect 13835 15668 13879 15706
rect 13761 15634 13879 15668
rect 13761 15600 13801 15634
rect 13835 15600 13879 15634
rect 13761 15566 13879 15600
rect 13761 15528 13801 15566
rect 13835 15528 13879 15566
rect 13761 15498 13879 15528
rect 13761 15456 13801 15498
rect 13835 15456 13879 15498
rect 13761 15430 13879 15456
rect 13761 15384 13801 15430
rect 13835 15384 13879 15430
rect 13761 15332 13879 15384
rect 1111 15291 13879 15332
rect 1111 15257 1290 15291
rect 1328 15257 1362 15291
rect 1396 15257 1430 15291
rect 1468 15257 1498 15291
rect 1540 15257 1566 15291
rect 1612 15257 1634 15291
rect 1684 15257 1702 15291
rect 1756 15257 1770 15291
rect 1828 15257 1838 15291
rect 1900 15257 1906 15291
rect 1972 15257 1974 15291
rect 2008 15257 2010 15291
rect 2076 15257 2082 15291
rect 2144 15257 2154 15291
rect 2212 15257 2226 15291
rect 2280 15257 2298 15291
rect 2348 15257 2370 15291
rect 2416 15257 2442 15291
rect 2484 15257 2514 15291
rect 2552 15257 2586 15291
rect 2620 15257 2654 15291
rect 2692 15257 2722 15291
rect 2764 15257 2790 15291
rect 2836 15257 2858 15291
rect 2908 15257 2926 15291
rect 2980 15257 2994 15291
rect 3052 15257 3062 15291
rect 3124 15257 3130 15291
rect 3196 15257 3198 15291
rect 3232 15257 3234 15291
rect 3300 15257 3306 15291
rect 3368 15257 3378 15291
rect 3436 15257 3450 15291
rect 3504 15257 3522 15291
rect 3572 15257 3594 15291
rect 3640 15257 3666 15291
rect 3708 15257 3738 15291
rect 3776 15257 3810 15291
rect 3844 15257 3878 15291
rect 3916 15257 3946 15291
rect 3988 15257 4014 15291
rect 4060 15257 4082 15291
rect 4132 15257 4150 15291
rect 4204 15257 4218 15291
rect 4276 15257 4286 15291
rect 4348 15257 4354 15291
rect 4420 15257 4422 15291
rect 4456 15257 4458 15291
rect 4524 15257 4530 15291
rect 4592 15257 4602 15291
rect 4660 15257 4674 15291
rect 4728 15257 4746 15291
rect 4796 15257 4818 15291
rect 4864 15257 4890 15291
rect 4932 15257 4962 15291
rect 5000 15257 5034 15291
rect 5068 15257 5102 15291
rect 5140 15257 5170 15291
rect 5212 15257 5238 15291
rect 5284 15257 5306 15291
rect 5356 15257 5374 15291
rect 5428 15257 5442 15291
rect 5500 15257 5510 15291
rect 5572 15257 5578 15291
rect 5644 15257 5646 15291
rect 5680 15257 5682 15291
rect 5748 15257 5754 15291
rect 5816 15257 5826 15291
rect 5884 15257 5898 15291
rect 5952 15257 5970 15291
rect 6020 15257 6042 15291
rect 6088 15257 6114 15291
rect 6156 15257 6186 15291
rect 6224 15257 6258 15291
rect 6292 15257 6326 15291
rect 6364 15257 6394 15291
rect 6436 15257 6462 15291
rect 6508 15257 6530 15291
rect 6580 15257 6598 15291
rect 6652 15257 6666 15291
rect 6724 15257 6734 15291
rect 6796 15257 6802 15291
rect 6868 15257 6870 15291
rect 6904 15257 6906 15291
rect 6972 15257 6978 15291
rect 7040 15257 7050 15291
rect 7108 15257 7122 15291
rect 7176 15257 7194 15291
rect 7244 15257 7266 15291
rect 7312 15257 7338 15291
rect 7380 15257 7410 15291
rect 7448 15257 7482 15291
rect 7516 15257 7550 15291
rect 7588 15257 7618 15291
rect 7660 15257 7686 15291
rect 7732 15257 7754 15291
rect 7804 15257 7822 15291
rect 7876 15257 7890 15291
rect 7948 15257 7958 15291
rect 8020 15257 8026 15291
rect 8092 15257 8094 15291
rect 8128 15257 8130 15291
rect 8196 15257 8202 15291
rect 8264 15257 8274 15291
rect 8332 15257 8346 15291
rect 8400 15257 8418 15291
rect 8468 15257 8490 15291
rect 8536 15257 8562 15291
rect 8604 15257 8634 15291
rect 8672 15257 8706 15291
rect 8740 15257 8774 15291
rect 8812 15257 8842 15291
rect 8884 15257 8910 15291
rect 8956 15257 8978 15291
rect 9028 15257 9046 15291
rect 9100 15257 9114 15291
rect 9172 15257 9182 15291
rect 9244 15257 9250 15291
rect 9316 15257 9318 15291
rect 9352 15257 9354 15291
rect 9420 15257 9426 15291
rect 9488 15257 9498 15291
rect 9556 15257 9570 15291
rect 9624 15257 9642 15291
rect 9692 15257 9714 15291
rect 9760 15257 9786 15291
rect 9828 15257 9858 15291
rect 9896 15257 9930 15291
rect 9964 15257 9998 15291
rect 10036 15257 10066 15291
rect 10108 15257 10134 15291
rect 10180 15257 10202 15291
rect 10252 15257 10270 15291
rect 10324 15257 10338 15291
rect 10396 15257 10406 15291
rect 10468 15257 10474 15291
rect 10540 15257 10542 15291
rect 10576 15257 10578 15291
rect 10644 15257 10650 15291
rect 10712 15257 10722 15291
rect 10780 15257 10794 15291
rect 10848 15257 10866 15291
rect 10916 15257 10938 15291
rect 10984 15257 11010 15291
rect 11052 15257 11082 15291
rect 11120 15257 11154 15291
rect 11188 15257 11222 15291
rect 11260 15257 11290 15291
rect 11332 15257 11358 15291
rect 11404 15257 11426 15291
rect 11476 15257 11494 15291
rect 11548 15257 11562 15291
rect 11620 15257 11630 15291
rect 11692 15257 11698 15291
rect 11764 15257 11766 15291
rect 11800 15257 11802 15291
rect 11868 15257 11874 15291
rect 11936 15257 11946 15291
rect 12004 15257 12018 15291
rect 12072 15257 12090 15291
rect 12140 15257 12162 15291
rect 12208 15257 12234 15291
rect 12276 15257 12306 15291
rect 12344 15257 12378 15291
rect 12412 15257 12446 15291
rect 12484 15257 12514 15291
rect 12556 15257 12582 15291
rect 12628 15257 12650 15291
rect 12700 15257 12718 15291
rect 12772 15257 12786 15291
rect 12844 15257 12854 15291
rect 12916 15257 12922 15291
rect 12988 15257 12990 15291
rect 13024 15257 13026 15291
rect 13092 15257 13098 15291
rect 13160 15257 13170 15291
rect 13228 15257 13242 15291
rect 13296 15257 13314 15291
rect 13364 15257 13386 15291
rect 13432 15257 13458 15291
rect 13500 15257 13530 15291
rect 13568 15257 13602 15291
rect 13636 15257 13670 15291
rect 13708 15257 13879 15291
rect 1111 15214 13879 15257
rect 13960 34720 14114 34754
rect 14148 34737 14289 34754
rect 14323 34737 14353 34771
rect 14148 34720 14353 34737
rect 13960 34703 14353 34720
rect 13960 34682 14289 34703
rect 13960 34648 14114 34682
rect 14148 34669 14289 34682
rect 14323 34669 14353 34703
rect 14148 34648 14353 34669
rect 13960 34635 14353 34648
rect 13960 34610 14289 34635
rect 13960 34576 14114 34610
rect 14148 34601 14289 34610
rect 14323 34601 14353 34635
rect 14148 34576 14353 34601
rect 13960 34567 14353 34576
rect 13960 34538 14289 34567
rect 13960 34504 14114 34538
rect 14148 34533 14289 34538
rect 14323 34533 14353 34567
rect 14148 34504 14353 34533
rect 13960 34499 14353 34504
rect 13960 34466 14289 34499
rect 13960 34432 14114 34466
rect 14148 34465 14289 34466
rect 14323 34465 14353 34499
rect 14148 34432 14353 34465
rect 13960 34431 14353 34432
rect 13960 34397 14289 34431
rect 14323 34397 14353 34431
rect 13960 34394 14353 34397
rect 13960 34360 14114 34394
rect 14148 34363 14353 34394
rect 14148 34360 14289 34363
rect 13960 34329 14289 34360
rect 14323 34329 14353 34363
rect 13960 34322 14353 34329
rect 13960 34288 14114 34322
rect 14148 34295 14353 34322
rect 14148 34288 14289 34295
rect 13960 34261 14289 34288
rect 14323 34261 14353 34295
rect 13960 34250 14353 34261
rect 13960 34216 14114 34250
rect 14148 34227 14353 34250
rect 14148 34216 14289 34227
rect 13960 34193 14289 34216
rect 14323 34193 14353 34227
rect 13960 34178 14353 34193
rect 13960 34144 14114 34178
rect 14148 34159 14353 34178
rect 14148 34144 14289 34159
rect 13960 34125 14289 34144
rect 14323 34125 14353 34159
rect 13960 34106 14353 34125
rect 13960 34072 14114 34106
rect 14148 34091 14353 34106
rect 14148 34072 14289 34091
rect 13960 34057 14289 34072
rect 14323 34057 14353 34091
rect 13960 34034 14353 34057
rect 13960 34000 14114 34034
rect 14148 34023 14353 34034
rect 14148 34000 14289 34023
rect 13960 33989 14289 34000
rect 14323 33989 14353 34023
rect 13960 33962 14353 33989
rect 13960 33928 14114 33962
rect 14148 33955 14353 33962
rect 14148 33928 14289 33955
rect 13960 33921 14289 33928
rect 14323 33921 14353 33955
rect 13960 33890 14353 33921
rect 13960 33856 14114 33890
rect 14148 33887 14353 33890
rect 14148 33856 14289 33887
rect 13960 33853 14289 33856
rect 14323 33853 14353 33887
rect 13960 33819 14353 33853
rect 13960 33818 14289 33819
rect 13960 33784 14114 33818
rect 14148 33785 14289 33818
rect 14323 33785 14353 33819
rect 14148 33784 14353 33785
rect 13960 33751 14353 33784
rect 13960 33746 14289 33751
rect 13960 33712 14114 33746
rect 14148 33717 14289 33746
rect 14323 33717 14353 33751
rect 14148 33712 14353 33717
rect 13960 33683 14353 33712
rect 13960 33674 14289 33683
rect 13960 33640 14114 33674
rect 14148 33649 14289 33674
rect 14323 33649 14353 33683
rect 14148 33640 14353 33649
rect 13960 33615 14353 33640
rect 13960 33602 14289 33615
rect 13960 33568 14114 33602
rect 14148 33581 14289 33602
rect 14323 33581 14353 33615
rect 14148 33568 14353 33581
rect 13960 33547 14353 33568
rect 13960 33530 14289 33547
rect 13960 33496 14114 33530
rect 14148 33513 14289 33530
rect 14323 33513 14353 33547
rect 14148 33496 14353 33513
rect 13960 33479 14353 33496
rect 13960 33458 14289 33479
rect 13960 33424 14114 33458
rect 14148 33445 14289 33458
rect 14323 33445 14353 33479
rect 14148 33424 14353 33445
rect 13960 33411 14353 33424
rect 13960 33386 14289 33411
rect 13960 33352 14114 33386
rect 14148 33377 14289 33386
rect 14323 33377 14353 33411
rect 14148 33352 14353 33377
rect 13960 33343 14353 33352
rect 13960 33314 14289 33343
rect 13960 33280 14114 33314
rect 14148 33309 14289 33314
rect 14323 33309 14353 33343
rect 14148 33280 14353 33309
rect 13960 33275 14353 33280
rect 13960 33242 14289 33275
rect 13960 33208 14114 33242
rect 14148 33241 14289 33242
rect 14323 33241 14353 33275
rect 14148 33208 14353 33241
rect 13960 33207 14353 33208
rect 13960 33173 14289 33207
rect 14323 33173 14353 33207
rect 13960 33170 14353 33173
rect 13960 33136 14114 33170
rect 14148 33139 14353 33170
rect 14148 33136 14289 33139
rect 13960 33105 14289 33136
rect 14323 33105 14353 33139
rect 13960 33098 14353 33105
rect 13960 33064 14114 33098
rect 14148 33071 14353 33098
rect 14148 33064 14289 33071
rect 13960 33037 14289 33064
rect 14323 33037 14353 33071
rect 13960 33026 14353 33037
rect 13960 32992 14114 33026
rect 14148 33003 14353 33026
rect 14148 32992 14289 33003
rect 13960 32969 14289 32992
rect 14323 32969 14353 33003
rect 13960 32954 14353 32969
rect 13960 32920 14114 32954
rect 14148 32935 14353 32954
rect 14148 32920 14289 32935
rect 13960 32901 14289 32920
rect 14323 32901 14353 32935
rect 13960 32882 14353 32901
rect 13960 32848 14114 32882
rect 14148 32867 14353 32882
rect 14148 32848 14289 32867
rect 13960 32833 14289 32848
rect 14323 32833 14353 32867
rect 13960 32810 14353 32833
rect 13960 32776 14114 32810
rect 14148 32799 14353 32810
rect 14148 32776 14289 32799
rect 13960 32765 14289 32776
rect 14323 32765 14353 32799
rect 13960 32738 14353 32765
rect 13960 32704 14114 32738
rect 14148 32731 14353 32738
rect 14148 32704 14289 32731
rect 13960 32697 14289 32704
rect 14323 32697 14353 32731
rect 13960 32666 14353 32697
rect 13960 32632 14114 32666
rect 14148 32663 14353 32666
rect 14148 32632 14289 32663
rect 13960 32629 14289 32632
rect 14323 32629 14353 32663
rect 13960 32595 14353 32629
rect 13960 32594 14289 32595
rect 13960 32560 14114 32594
rect 14148 32561 14289 32594
rect 14323 32561 14353 32595
rect 14148 32560 14353 32561
rect 13960 32527 14353 32560
rect 13960 32522 14289 32527
rect 13960 32488 14114 32522
rect 14148 32493 14289 32522
rect 14323 32493 14353 32527
rect 14148 32488 14353 32493
rect 13960 32459 14353 32488
rect 13960 32450 14289 32459
rect 13960 32416 14114 32450
rect 14148 32425 14289 32450
rect 14323 32425 14353 32459
rect 14148 32416 14353 32425
rect 13960 32391 14353 32416
rect 13960 32378 14289 32391
rect 13960 32344 14114 32378
rect 14148 32357 14289 32378
rect 14323 32357 14353 32391
rect 14148 32344 14353 32357
rect 13960 32323 14353 32344
rect 13960 32306 14289 32323
rect 13960 32272 14114 32306
rect 14148 32289 14289 32306
rect 14323 32289 14353 32323
rect 14148 32272 14353 32289
rect 13960 32255 14353 32272
rect 13960 32234 14289 32255
rect 13960 32200 14114 32234
rect 14148 32221 14289 32234
rect 14323 32221 14353 32255
rect 14148 32200 14353 32221
rect 13960 32187 14353 32200
rect 13960 32162 14289 32187
rect 13960 32128 14114 32162
rect 14148 32153 14289 32162
rect 14323 32153 14353 32187
rect 14148 32128 14353 32153
rect 13960 32119 14353 32128
rect 13960 32090 14289 32119
rect 13960 32056 14114 32090
rect 14148 32085 14289 32090
rect 14323 32085 14353 32119
rect 14148 32056 14353 32085
rect 13960 32051 14353 32056
rect 13960 32018 14289 32051
rect 13960 31984 14114 32018
rect 14148 32017 14289 32018
rect 14323 32017 14353 32051
rect 14148 31984 14353 32017
rect 13960 31983 14353 31984
rect 13960 31949 14289 31983
rect 14323 31949 14353 31983
rect 13960 31946 14353 31949
rect 13960 31912 14114 31946
rect 14148 31915 14353 31946
rect 14148 31912 14289 31915
rect 13960 31881 14289 31912
rect 14323 31881 14353 31915
rect 13960 31874 14353 31881
rect 13960 31840 14114 31874
rect 14148 31847 14353 31874
rect 14148 31840 14289 31847
rect 13960 31813 14289 31840
rect 14323 31813 14353 31847
rect 13960 31802 14353 31813
rect 13960 31768 14114 31802
rect 14148 31779 14353 31802
rect 14148 31768 14289 31779
rect 13960 31745 14289 31768
rect 14323 31745 14353 31779
rect 13960 31730 14353 31745
rect 13960 31696 14114 31730
rect 14148 31711 14353 31730
rect 14148 31696 14289 31711
rect 13960 31677 14289 31696
rect 14323 31677 14353 31711
rect 13960 31658 14353 31677
rect 13960 31624 14114 31658
rect 14148 31643 14353 31658
rect 14148 31624 14289 31643
rect 13960 31609 14289 31624
rect 14323 31609 14353 31643
rect 13960 31586 14353 31609
rect 13960 31552 14114 31586
rect 14148 31575 14353 31586
rect 14148 31552 14289 31575
rect 13960 31541 14289 31552
rect 14323 31541 14353 31575
rect 13960 31514 14353 31541
rect 13960 31480 14114 31514
rect 14148 31507 14353 31514
rect 14148 31480 14289 31507
rect 13960 31473 14289 31480
rect 14323 31473 14353 31507
rect 13960 31442 14353 31473
rect 13960 31408 14114 31442
rect 14148 31439 14353 31442
rect 14148 31408 14289 31439
rect 13960 31405 14289 31408
rect 14323 31405 14353 31439
rect 13960 31371 14353 31405
rect 13960 31370 14289 31371
rect 13960 31336 14114 31370
rect 14148 31337 14289 31370
rect 14323 31337 14353 31371
rect 14148 31336 14353 31337
rect 13960 31303 14353 31336
rect 13960 31298 14289 31303
rect 13960 31264 14114 31298
rect 14148 31269 14289 31298
rect 14323 31269 14353 31303
rect 14148 31264 14353 31269
rect 13960 31235 14353 31264
rect 13960 31226 14289 31235
rect 13960 31192 14114 31226
rect 14148 31201 14289 31226
rect 14323 31201 14353 31235
rect 14148 31192 14353 31201
rect 13960 31167 14353 31192
rect 13960 31154 14289 31167
rect 13960 31120 14114 31154
rect 14148 31133 14289 31154
rect 14323 31133 14353 31167
rect 14148 31120 14353 31133
rect 13960 31099 14353 31120
rect 13960 31082 14289 31099
rect 13960 31048 14114 31082
rect 14148 31065 14289 31082
rect 14323 31065 14353 31099
rect 14148 31048 14353 31065
rect 13960 31031 14353 31048
rect 13960 31010 14289 31031
rect 13960 30976 14114 31010
rect 14148 30997 14289 31010
rect 14323 30997 14353 31031
rect 14148 30976 14353 30997
rect 13960 30963 14353 30976
rect 13960 30938 14289 30963
rect 13960 30904 14114 30938
rect 14148 30929 14289 30938
rect 14323 30929 14353 30963
rect 14148 30904 14353 30929
rect 13960 30895 14353 30904
rect 13960 30866 14289 30895
rect 13960 30832 14114 30866
rect 14148 30861 14289 30866
rect 14323 30861 14353 30895
rect 14148 30832 14353 30861
rect 13960 30827 14353 30832
rect 13960 30794 14289 30827
rect 13960 30760 14114 30794
rect 14148 30793 14289 30794
rect 14323 30793 14353 30827
rect 14148 30760 14353 30793
rect 13960 30759 14353 30760
rect 13960 30725 14289 30759
rect 14323 30725 14353 30759
rect 13960 30722 14353 30725
rect 13960 30688 14114 30722
rect 14148 30691 14353 30722
rect 14148 30688 14289 30691
rect 13960 30657 14289 30688
rect 14323 30657 14353 30691
rect 13960 30650 14353 30657
rect 13960 30616 14114 30650
rect 14148 30623 14353 30650
rect 14148 30616 14289 30623
rect 13960 30589 14289 30616
rect 14323 30589 14353 30623
rect 13960 30578 14353 30589
rect 13960 30544 14114 30578
rect 14148 30555 14353 30578
rect 14148 30544 14289 30555
rect 13960 30521 14289 30544
rect 14323 30521 14353 30555
rect 13960 30506 14353 30521
rect 13960 30472 14114 30506
rect 14148 30487 14353 30506
rect 14148 30472 14289 30487
rect 13960 30453 14289 30472
rect 14323 30453 14353 30487
rect 13960 30434 14353 30453
rect 13960 30400 14114 30434
rect 14148 30419 14353 30434
rect 14148 30400 14289 30419
rect 13960 30385 14289 30400
rect 14323 30385 14353 30419
rect 13960 30362 14353 30385
rect 13960 30328 14114 30362
rect 14148 30351 14353 30362
rect 14148 30328 14289 30351
rect 13960 30317 14289 30328
rect 14323 30317 14353 30351
rect 13960 30290 14353 30317
rect 13960 30256 14114 30290
rect 14148 30283 14353 30290
rect 14148 30256 14289 30283
rect 13960 30249 14289 30256
rect 14323 30249 14353 30283
rect 13960 30218 14353 30249
rect 13960 30184 14114 30218
rect 14148 30215 14353 30218
rect 14148 30184 14289 30215
rect 13960 30181 14289 30184
rect 14323 30181 14353 30215
rect 13960 30147 14353 30181
rect 13960 30146 14289 30147
rect 13960 30112 14114 30146
rect 14148 30113 14289 30146
rect 14323 30113 14353 30147
rect 14148 30112 14353 30113
rect 13960 30079 14353 30112
rect 13960 30074 14289 30079
rect 13960 30040 14114 30074
rect 14148 30045 14289 30074
rect 14323 30045 14353 30079
rect 14148 30040 14353 30045
rect 13960 30011 14353 30040
rect 13960 30002 14289 30011
rect 13960 29968 14114 30002
rect 14148 29977 14289 30002
rect 14323 29977 14353 30011
rect 14148 29968 14353 29977
rect 13960 29943 14353 29968
rect 13960 29930 14289 29943
rect 13960 29896 14114 29930
rect 14148 29909 14289 29930
rect 14323 29909 14353 29943
rect 14148 29896 14353 29909
rect 13960 29875 14353 29896
rect 13960 29858 14289 29875
rect 13960 29824 14114 29858
rect 14148 29841 14289 29858
rect 14323 29841 14353 29875
rect 14148 29824 14353 29841
rect 13960 29807 14353 29824
rect 13960 29786 14289 29807
rect 13960 29752 14114 29786
rect 14148 29773 14289 29786
rect 14323 29773 14353 29807
rect 14148 29752 14353 29773
rect 13960 29739 14353 29752
rect 13960 29714 14289 29739
rect 13960 29680 14114 29714
rect 14148 29705 14289 29714
rect 14323 29705 14353 29739
rect 14148 29680 14353 29705
rect 13960 29671 14353 29680
rect 13960 29642 14289 29671
rect 13960 29608 14114 29642
rect 14148 29637 14289 29642
rect 14323 29637 14353 29671
rect 14148 29608 14353 29637
rect 13960 29603 14353 29608
rect 13960 29570 14289 29603
rect 13960 29536 14114 29570
rect 14148 29569 14289 29570
rect 14323 29569 14353 29603
rect 14148 29536 14353 29569
rect 13960 29535 14353 29536
rect 13960 29501 14289 29535
rect 14323 29501 14353 29535
rect 13960 29498 14353 29501
rect 13960 29464 14114 29498
rect 14148 29467 14353 29498
rect 14148 29464 14289 29467
rect 13960 29433 14289 29464
rect 14323 29433 14353 29467
rect 13960 29426 14353 29433
rect 13960 29392 14114 29426
rect 14148 29399 14353 29426
rect 14148 29392 14289 29399
rect 13960 29365 14289 29392
rect 14323 29365 14353 29399
rect 13960 29354 14353 29365
rect 13960 29320 14114 29354
rect 14148 29331 14353 29354
rect 14148 29320 14289 29331
rect 13960 29297 14289 29320
rect 14323 29297 14353 29331
rect 13960 29282 14353 29297
rect 13960 29248 14114 29282
rect 14148 29263 14353 29282
rect 14148 29248 14289 29263
rect 13960 29229 14289 29248
rect 14323 29229 14353 29263
rect 13960 29210 14353 29229
rect 13960 29176 14114 29210
rect 14148 29195 14353 29210
rect 14148 29176 14289 29195
rect 13960 29161 14289 29176
rect 14323 29161 14353 29195
rect 13960 29138 14353 29161
rect 13960 29104 14114 29138
rect 14148 29127 14353 29138
rect 14148 29104 14289 29127
rect 13960 29093 14289 29104
rect 14323 29093 14353 29127
rect 13960 29066 14353 29093
rect 13960 29032 14114 29066
rect 14148 29059 14353 29066
rect 14148 29032 14289 29059
rect 13960 29025 14289 29032
rect 14323 29025 14353 29059
rect 13960 28994 14353 29025
rect 13960 28960 14114 28994
rect 14148 28991 14353 28994
rect 14148 28960 14289 28991
rect 13960 28957 14289 28960
rect 14323 28957 14353 28991
rect 13960 28923 14353 28957
rect 13960 28922 14289 28923
rect 13960 28888 14114 28922
rect 14148 28889 14289 28922
rect 14323 28889 14353 28923
rect 14148 28888 14353 28889
rect 13960 28855 14353 28888
rect 13960 28850 14289 28855
rect 13960 28816 14114 28850
rect 14148 28821 14289 28850
rect 14323 28821 14353 28855
rect 14148 28816 14353 28821
rect 13960 28787 14353 28816
rect 13960 28778 14289 28787
rect 13960 28744 14114 28778
rect 14148 28753 14289 28778
rect 14323 28753 14353 28787
rect 14148 28744 14353 28753
rect 13960 28719 14353 28744
rect 13960 28706 14289 28719
rect 13960 28672 14114 28706
rect 14148 28685 14289 28706
rect 14323 28685 14353 28719
rect 14148 28672 14353 28685
rect 13960 28651 14353 28672
rect 13960 28634 14289 28651
rect 13960 28600 14114 28634
rect 14148 28617 14289 28634
rect 14323 28617 14353 28651
rect 14148 28600 14353 28617
rect 13960 28583 14353 28600
rect 13960 28562 14289 28583
rect 13960 28528 14114 28562
rect 14148 28549 14289 28562
rect 14323 28549 14353 28583
rect 14148 28528 14353 28549
rect 13960 28515 14353 28528
rect 13960 28490 14289 28515
rect 13960 28456 14114 28490
rect 14148 28481 14289 28490
rect 14323 28481 14353 28515
rect 14148 28456 14353 28481
rect 13960 28447 14353 28456
rect 13960 28418 14289 28447
rect 13960 28384 14114 28418
rect 14148 28413 14289 28418
rect 14323 28413 14353 28447
rect 14148 28384 14353 28413
rect 13960 28379 14353 28384
rect 13960 28346 14289 28379
rect 13960 28312 14114 28346
rect 14148 28345 14289 28346
rect 14323 28345 14353 28379
rect 14148 28312 14353 28345
rect 13960 28311 14353 28312
rect 13960 28277 14289 28311
rect 14323 28277 14353 28311
rect 13960 28274 14353 28277
rect 13960 28240 14114 28274
rect 14148 28243 14353 28274
rect 14148 28240 14289 28243
rect 13960 28209 14289 28240
rect 14323 28209 14353 28243
rect 13960 28202 14353 28209
rect 13960 28168 14114 28202
rect 14148 28175 14353 28202
rect 14148 28168 14289 28175
rect 13960 28141 14289 28168
rect 14323 28141 14353 28175
rect 13960 28130 14353 28141
rect 13960 28096 14114 28130
rect 14148 28107 14353 28130
rect 14148 28096 14289 28107
rect 13960 28073 14289 28096
rect 14323 28073 14353 28107
rect 13960 28058 14353 28073
rect 13960 28024 14114 28058
rect 14148 28039 14353 28058
rect 14148 28024 14289 28039
rect 13960 28005 14289 28024
rect 14323 28005 14353 28039
rect 13960 27986 14353 28005
rect 13960 27952 14114 27986
rect 14148 27971 14353 27986
rect 14148 27952 14289 27971
rect 13960 27937 14289 27952
rect 14323 27937 14353 27971
rect 13960 27914 14353 27937
rect 13960 27880 14114 27914
rect 14148 27903 14353 27914
rect 14148 27880 14289 27903
rect 13960 27869 14289 27880
rect 14323 27869 14353 27903
rect 13960 27842 14353 27869
rect 13960 27808 14114 27842
rect 14148 27835 14353 27842
rect 14148 27808 14289 27835
rect 13960 27801 14289 27808
rect 14323 27801 14353 27835
rect 13960 27770 14353 27801
rect 13960 27736 14114 27770
rect 14148 27767 14353 27770
rect 14148 27736 14289 27767
rect 13960 27733 14289 27736
rect 14323 27733 14353 27767
rect 13960 27699 14353 27733
rect 13960 27698 14289 27699
rect 13960 27664 14114 27698
rect 14148 27665 14289 27698
rect 14323 27665 14353 27699
rect 14148 27664 14353 27665
rect 13960 27631 14353 27664
rect 13960 27626 14289 27631
rect 13960 27592 14114 27626
rect 14148 27597 14289 27626
rect 14323 27597 14353 27631
rect 14148 27592 14353 27597
rect 13960 27563 14353 27592
rect 13960 27554 14289 27563
rect 13960 27520 14114 27554
rect 14148 27529 14289 27554
rect 14323 27529 14353 27563
rect 14148 27520 14353 27529
rect 13960 27495 14353 27520
rect 13960 27482 14289 27495
rect 13960 27448 14114 27482
rect 14148 27461 14289 27482
rect 14323 27461 14353 27495
rect 14148 27448 14353 27461
rect 13960 27427 14353 27448
rect 13960 27410 14289 27427
rect 13960 27376 14114 27410
rect 14148 27393 14289 27410
rect 14323 27393 14353 27427
rect 14148 27376 14353 27393
rect 13960 27359 14353 27376
rect 13960 27338 14289 27359
rect 13960 27304 14114 27338
rect 14148 27325 14289 27338
rect 14323 27325 14353 27359
rect 14148 27304 14353 27325
rect 13960 27291 14353 27304
rect 13960 27266 14289 27291
rect 13960 27232 14114 27266
rect 14148 27257 14289 27266
rect 14323 27257 14353 27291
rect 14148 27232 14353 27257
rect 13960 27223 14353 27232
rect 13960 27194 14289 27223
rect 13960 27160 14114 27194
rect 14148 27189 14289 27194
rect 14323 27189 14353 27223
rect 14148 27160 14353 27189
rect 13960 27155 14353 27160
rect 13960 27122 14289 27155
rect 13960 27088 14114 27122
rect 14148 27121 14289 27122
rect 14323 27121 14353 27155
rect 14148 27088 14353 27121
rect 13960 27087 14353 27088
rect 13960 27053 14289 27087
rect 14323 27053 14353 27087
rect 13960 27050 14353 27053
rect 13960 27016 14114 27050
rect 14148 27019 14353 27050
rect 14148 27016 14289 27019
rect 13960 26985 14289 27016
rect 14323 26985 14353 27019
rect 13960 26978 14353 26985
rect 13960 26944 14114 26978
rect 14148 26951 14353 26978
rect 14148 26944 14289 26951
rect 13960 26917 14289 26944
rect 14323 26917 14353 26951
rect 13960 26906 14353 26917
rect 13960 26872 14114 26906
rect 14148 26883 14353 26906
rect 14148 26872 14289 26883
rect 13960 26849 14289 26872
rect 14323 26849 14353 26883
rect 13960 26834 14353 26849
rect 13960 26800 14114 26834
rect 14148 26815 14353 26834
rect 14148 26800 14289 26815
rect 13960 26781 14289 26800
rect 14323 26781 14353 26815
rect 13960 26762 14353 26781
rect 13960 26728 14114 26762
rect 14148 26747 14353 26762
rect 14148 26728 14289 26747
rect 13960 26713 14289 26728
rect 14323 26713 14353 26747
rect 13960 26690 14353 26713
rect 13960 26656 14114 26690
rect 14148 26679 14353 26690
rect 14148 26656 14289 26679
rect 13960 26645 14289 26656
rect 14323 26645 14353 26679
rect 13960 26618 14353 26645
rect 13960 26584 14114 26618
rect 14148 26611 14353 26618
rect 14148 26584 14289 26611
rect 13960 26577 14289 26584
rect 14323 26577 14353 26611
rect 13960 26546 14353 26577
rect 13960 26512 14114 26546
rect 14148 26543 14353 26546
rect 14148 26512 14289 26543
rect 13960 26509 14289 26512
rect 14323 26509 14353 26543
rect 13960 26475 14353 26509
rect 13960 26474 14289 26475
rect 13960 26440 14114 26474
rect 14148 26441 14289 26474
rect 14323 26441 14353 26475
rect 14148 26440 14353 26441
rect 13960 26407 14353 26440
rect 13960 26402 14289 26407
rect 13960 26368 14114 26402
rect 14148 26373 14289 26402
rect 14323 26373 14353 26407
rect 14148 26368 14353 26373
rect 13960 26339 14353 26368
rect 13960 26330 14289 26339
rect 13960 26296 14114 26330
rect 14148 26305 14289 26330
rect 14323 26305 14353 26339
rect 14148 26296 14353 26305
rect 13960 26271 14353 26296
rect 13960 26258 14289 26271
rect 13960 26224 14114 26258
rect 14148 26237 14289 26258
rect 14323 26237 14353 26271
rect 14148 26224 14353 26237
rect 13960 26203 14353 26224
rect 13960 26186 14289 26203
rect 13960 26152 14114 26186
rect 14148 26169 14289 26186
rect 14323 26169 14353 26203
rect 14148 26152 14353 26169
rect 13960 26135 14353 26152
rect 13960 26114 14289 26135
rect 13960 26080 14114 26114
rect 14148 26101 14289 26114
rect 14323 26101 14353 26135
rect 14148 26080 14353 26101
rect 13960 26067 14353 26080
rect 13960 26042 14289 26067
rect 13960 26008 14114 26042
rect 14148 26033 14289 26042
rect 14323 26033 14353 26067
rect 14148 26008 14353 26033
rect 13960 25999 14353 26008
rect 13960 25970 14289 25999
rect 13960 25936 14114 25970
rect 14148 25965 14289 25970
rect 14323 25965 14353 25999
rect 14148 25936 14353 25965
rect 13960 25931 14353 25936
rect 13960 25898 14289 25931
rect 13960 25864 14114 25898
rect 14148 25897 14289 25898
rect 14323 25897 14353 25931
rect 14148 25864 14353 25897
rect 13960 25863 14353 25864
rect 13960 25829 14289 25863
rect 14323 25829 14353 25863
rect 13960 25826 14353 25829
rect 13960 25792 14114 25826
rect 14148 25795 14353 25826
rect 14148 25792 14289 25795
rect 13960 25761 14289 25792
rect 14323 25761 14353 25795
rect 13960 25754 14353 25761
rect 13960 25720 14114 25754
rect 14148 25727 14353 25754
rect 14148 25720 14289 25727
rect 13960 25693 14289 25720
rect 14323 25693 14353 25727
rect 13960 25682 14353 25693
rect 13960 25648 14114 25682
rect 14148 25659 14353 25682
rect 14148 25648 14289 25659
rect 13960 25625 14289 25648
rect 14323 25625 14353 25659
rect 13960 25610 14353 25625
rect 13960 25576 14114 25610
rect 14148 25591 14353 25610
rect 14148 25576 14289 25591
rect 13960 25557 14289 25576
rect 14323 25557 14353 25591
rect 13960 25538 14353 25557
rect 13960 25504 14114 25538
rect 14148 25523 14353 25538
rect 14148 25504 14289 25523
rect 13960 25489 14289 25504
rect 14323 25489 14353 25523
rect 13960 25466 14353 25489
rect 13960 25432 14114 25466
rect 14148 25455 14353 25466
rect 14148 25432 14289 25455
rect 13960 25421 14289 25432
rect 14323 25421 14353 25455
rect 13960 25394 14353 25421
rect 13960 25360 14114 25394
rect 14148 25387 14353 25394
rect 14148 25360 14289 25387
rect 13960 25353 14289 25360
rect 14323 25353 14353 25387
rect 13960 25322 14353 25353
rect 13960 25288 14114 25322
rect 14148 25319 14353 25322
rect 14148 25288 14289 25319
rect 13960 25285 14289 25288
rect 14323 25285 14353 25319
rect 13960 25251 14353 25285
rect 13960 25250 14289 25251
rect 13960 25216 14114 25250
rect 14148 25217 14289 25250
rect 14323 25217 14353 25251
rect 14148 25216 14353 25217
rect 13960 25183 14353 25216
rect 13960 25178 14289 25183
rect 13960 25144 14114 25178
rect 14148 25149 14289 25178
rect 14323 25149 14353 25183
rect 14148 25144 14353 25149
rect 13960 25115 14353 25144
rect 13960 25106 14289 25115
rect 13960 25072 14114 25106
rect 14148 25081 14289 25106
rect 14323 25081 14353 25115
rect 14148 25072 14353 25081
rect 13960 25047 14353 25072
rect 13960 25034 14289 25047
rect 13960 25000 14114 25034
rect 14148 25013 14289 25034
rect 14323 25013 14353 25047
rect 14148 25000 14353 25013
rect 13960 24979 14353 25000
rect 13960 24962 14289 24979
rect 13960 24928 14114 24962
rect 14148 24945 14289 24962
rect 14323 24945 14353 24979
rect 14148 24928 14353 24945
rect 13960 24911 14353 24928
rect 13960 24890 14289 24911
rect 13960 24856 14114 24890
rect 14148 24877 14289 24890
rect 14323 24877 14353 24911
rect 14148 24856 14353 24877
rect 13960 24843 14353 24856
rect 13960 24818 14289 24843
rect 13960 24784 14114 24818
rect 14148 24809 14289 24818
rect 14323 24809 14353 24843
rect 14148 24784 14353 24809
rect 13960 24775 14353 24784
rect 13960 24746 14289 24775
rect 13960 24712 14114 24746
rect 14148 24741 14289 24746
rect 14323 24741 14353 24775
rect 14148 24712 14353 24741
rect 13960 24707 14353 24712
rect 13960 24674 14289 24707
rect 13960 24640 14114 24674
rect 14148 24673 14289 24674
rect 14323 24673 14353 24707
rect 14148 24640 14353 24673
rect 13960 24639 14353 24640
rect 13960 24605 14289 24639
rect 14323 24605 14353 24639
rect 13960 24602 14353 24605
rect 13960 24568 14114 24602
rect 14148 24571 14353 24602
rect 14148 24568 14289 24571
rect 13960 24537 14289 24568
rect 14323 24537 14353 24571
rect 13960 24530 14353 24537
rect 13960 24496 14114 24530
rect 14148 24503 14353 24530
rect 14148 24496 14289 24503
rect 13960 24469 14289 24496
rect 14323 24469 14353 24503
rect 13960 24458 14353 24469
rect 13960 24424 14114 24458
rect 14148 24435 14353 24458
rect 14148 24424 14289 24435
rect 13960 24401 14289 24424
rect 14323 24401 14353 24435
rect 13960 24386 14353 24401
rect 13960 24352 14114 24386
rect 14148 24367 14353 24386
rect 14148 24352 14289 24367
rect 13960 24333 14289 24352
rect 14323 24333 14353 24367
rect 13960 24314 14353 24333
rect 13960 24280 14114 24314
rect 14148 24299 14353 24314
rect 14148 24280 14289 24299
rect 13960 24265 14289 24280
rect 14323 24265 14353 24299
rect 13960 24242 14353 24265
rect 13960 24208 14114 24242
rect 14148 24231 14353 24242
rect 14148 24208 14289 24231
rect 13960 24197 14289 24208
rect 14323 24197 14353 24231
rect 13960 24170 14353 24197
rect 13960 24136 14114 24170
rect 14148 24163 14353 24170
rect 14148 24136 14289 24163
rect 13960 24129 14289 24136
rect 14323 24129 14353 24163
rect 13960 24098 14353 24129
rect 13960 24064 14114 24098
rect 14148 24095 14353 24098
rect 14148 24064 14289 24095
rect 13960 24061 14289 24064
rect 14323 24061 14353 24095
rect 13960 24027 14353 24061
rect 13960 24026 14289 24027
rect 13960 23992 14114 24026
rect 14148 23993 14289 24026
rect 14323 23993 14353 24027
rect 14148 23992 14353 23993
rect 13960 23959 14353 23992
rect 13960 23954 14289 23959
rect 13960 23920 14114 23954
rect 14148 23925 14289 23954
rect 14323 23925 14353 23959
rect 14148 23920 14353 23925
rect 13960 23891 14353 23920
rect 13960 23882 14289 23891
rect 13960 23848 14114 23882
rect 14148 23857 14289 23882
rect 14323 23857 14353 23891
rect 14148 23848 14353 23857
rect 13960 23823 14353 23848
rect 13960 23810 14289 23823
rect 13960 23776 14114 23810
rect 14148 23789 14289 23810
rect 14323 23789 14353 23823
rect 14148 23776 14353 23789
rect 13960 23755 14353 23776
rect 13960 23738 14289 23755
rect 13960 23704 14114 23738
rect 14148 23721 14289 23738
rect 14323 23721 14353 23755
rect 14148 23704 14353 23721
rect 13960 23687 14353 23704
rect 13960 23666 14289 23687
rect 13960 23632 14114 23666
rect 14148 23653 14289 23666
rect 14323 23653 14353 23687
rect 14148 23632 14353 23653
rect 13960 23619 14353 23632
rect 13960 23594 14289 23619
rect 13960 23560 14114 23594
rect 14148 23585 14289 23594
rect 14323 23585 14353 23619
rect 14148 23560 14353 23585
rect 13960 23551 14353 23560
rect 13960 23522 14289 23551
rect 13960 23488 14114 23522
rect 14148 23517 14289 23522
rect 14323 23517 14353 23551
rect 14148 23488 14353 23517
rect 13960 23483 14353 23488
rect 13960 23450 14289 23483
rect 13960 23416 14114 23450
rect 14148 23449 14289 23450
rect 14323 23449 14353 23483
rect 14148 23416 14353 23449
rect 13960 23415 14353 23416
rect 13960 23381 14289 23415
rect 14323 23381 14353 23415
rect 13960 23378 14353 23381
rect 13960 23344 14114 23378
rect 14148 23347 14353 23378
rect 14148 23344 14289 23347
rect 13960 23313 14289 23344
rect 14323 23313 14353 23347
rect 13960 23306 14353 23313
rect 13960 23272 14114 23306
rect 14148 23279 14353 23306
rect 14148 23272 14289 23279
rect 13960 23245 14289 23272
rect 14323 23245 14353 23279
rect 13960 23234 14353 23245
rect 13960 23200 14114 23234
rect 14148 23211 14353 23234
rect 14148 23200 14289 23211
rect 13960 23177 14289 23200
rect 14323 23177 14353 23211
rect 13960 23162 14353 23177
rect 13960 23128 14114 23162
rect 14148 23143 14353 23162
rect 14148 23128 14289 23143
rect 13960 23109 14289 23128
rect 14323 23109 14353 23143
rect 13960 23090 14353 23109
rect 13960 23056 14114 23090
rect 14148 23075 14353 23090
rect 14148 23056 14289 23075
rect 13960 23041 14289 23056
rect 14323 23041 14353 23075
rect 13960 23018 14353 23041
rect 13960 22984 14114 23018
rect 14148 23007 14353 23018
rect 14148 22984 14289 23007
rect 13960 22973 14289 22984
rect 14323 22973 14353 23007
rect 13960 22946 14353 22973
rect 13960 22912 14114 22946
rect 14148 22939 14353 22946
rect 14148 22912 14289 22939
rect 13960 22905 14289 22912
rect 14323 22905 14353 22939
rect 13960 22874 14353 22905
rect 13960 22840 14114 22874
rect 14148 22871 14353 22874
rect 14148 22840 14289 22871
rect 13960 22837 14289 22840
rect 14323 22837 14353 22871
rect 13960 22803 14353 22837
rect 13960 22802 14289 22803
rect 13960 22768 14114 22802
rect 14148 22769 14289 22802
rect 14323 22769 14353 22803
rect 14148 22768 14353 22769
rect 13960 22735 14353 22768
rect 13960 22730 14289 22735
rect 13960 22696 14114 22730
rect 14148 22701 14289 22730
rect 14323 22701 14353 22735
rect 14148 22696 14353 22701
rect 13960 22667 14353 22696
rect 13960 22658 14289 22667
rect 13960 22624 14114 22658
rect 14148 22633 14289 22658
rect 14323 22633 14353 22667
rect 14148 22624 14353 22633
rect 13960 22599 14353 22624
rect 13960 22586 14289 22599
rect 13960 22552 14114 22586
rect 14148 22565 14289 22586
rect 14323 22565 14353 22599
rect 14148 22552 14353 22565
rect 13960 22531 14353 22552
rect 13960 22514 14289 22531
rect 13960 22480 14114 22514
rect 14148 22497 14289 22514
rect 14323 22497 14353 22531
rect 14148 22480 14353 22497
rect 13960 22463 14353 22480
rect 13960 22442 14289 22463
rect 13960 22408 14114 22442
rect 14148 22429 14289 22442
rect 14323 22429 14353 22463
rect 14148 22408 14353 22429
rect 13960 22395 14353 22408
rect 13960 22370 14289 22395
rect 13960 22336 14114 22370
rect 14148 22361 14289 22370
rect 14323 22361 14353 22395
rect 14148 22336 14353 22361
rect 13960 22327 14353 22336
rect 13960 22298 14289 22327
rect 13960 22264 14114 22298
rect 14148 22293 14289 22298
rect 14323 22293 14353 22327
rect 14148 22264 14353 22293
rect 13960 22259 14353 22264
rect 13960 22226 14289 22259
rect 13960 22192 14114 22226
rect 14148 22225 14289 22226
rect 14323 22225 14353 22259
rect 14148 22192 14353 22225
rect 13960 22191 14353 22192
rect 13960 22157 14289 22191
rect 14323 22157 14353 22191
rect 13960 22154 14353 22157
rect 13960 22120 14114 22154
rect 14148 22123 14353 22154
rect 14148 22120 14289 22123
rect 13960 22089 14289 22120
rect 14323 22089 14353 22123
rect 13960 22082 14353 22089
rect 13960 22048 14114 22082
rect 14148 22055 14353 22082
rect 14148 22048 14289 22055
rect 13960 22021 14289 22048
rect 14323 22021 14353 22055
rect 13960 22010 14353 22021
rect 13960 21976 14114 22010
rect 14148 21987 14353 22010
rect 14148 21976 14289 21987
rect 13960 21953 14289 21976
rect 14323 21953 14353 21987
rect 13960 21938 14353 21953
rect 13960 21904 14114 21938
rect 14148 21919 14353 21938
rect 14148 21904 14289 21919
rect 13960 21885 14289 21904
rect 14323 21885 14353 21919
rect 13960 21866 14353 21885
rect 13960 21832 14114 21866
rect 14148 21851 14353 21866
rect 14148 21832 14289 21851
rect 13960 21817 14289 21832
rect 14323 21817 14353 21851
rect 13960 21794 14353 21817
rect 13960 21760 14114 21794
rect 14148 21783 14353 21794
rect 14148 21760 14289 21783
rect 13960 21749 14289 21760
rect 14323 21749 14353 21783
rect 13960 21722 14353 21749
rect 13960 21688 14114 21722
rect 14148 21715 14353 21722
rect 14148 21688 14289 21715
rect 13960 21681 14289 21688
rect 14323 21681 14353 21715
rect 13960 21650 14353 21681
rect 13960 21616 14114 21650
rect 14148 21647 14353 21650
rect 14148 21616 14289 21647
rect 13960 21613 14289 21616
rect 14323 21613 14353 21647
rect 13960 21579 14353 21613
rect 13960 21578 14289 21579
rect 13960 21544 14114 21578
rect 14148 21545 14289 21578
rect 14323 21545 14353 21579
rect 14148 21544 14353 21545
rect 13960 21511 14353 21544
rect 13960 21506 14289 21511
rect 13960 21472 14114 21506
rect 14148 21477 14289 21506
rect 14323 21477 14353 21511
rect 14148 21472 14353 21477
rect 13960 21443 14353 21472
rect 13960 21434 14289 21443
rect 13960 21400 14114 21434
rect 14148 21409 14289 21434
rect 14323 21409 14353 21443
rect 14148 21400 14353 21409
rect 13960 21375 14353 21400
rect 13960 21362 14289 21375
rect 13960 21328 14114 21362
rect 14148 21341 14289 21362
rect 14323 21341 14353 21375
rect 14148 21328 14353 21341
rect 13960 21307 14353 21328
rect 13960 21290 14289 21307
rect 13960 21256 14114 21290
rect 14148 21273 14289 21290
rect 14323 21273 14353 21307
rect 14148 21256 14353 21273
rect 13960 21239 14353 21256
rect 13960 21218 14289 21239
rect 13960 21184 14114 21218
rect 14148 21205 14289 21218
rect 14323 21205 14353 21239
rect 14148 21184 14353 21205
rect 13960 21171 14353 21184
rect 13960 21146 14289 21171
rect 13960 21112 14114 21146
rect 14148 21137 14289 21146
rect 14323 21137 14353 21171
rect 14148 21112 14353 21137
rect 13960 21103 14353 21112
rect 13960 21074 14289 21103
rect 13960 21040 14114 21074
rect 14148 21069 14289 21074
rect 14323 21069 14353 21103
rect 14148 21040 14353 21069
rect 13960 21035 14353 21040
rect 13960 21002 14289 21035
rect 13960 20968 14114 21002
rect 14148 21001 14289 21002
rect 14323 21001 14353 21035
rect 14148 20968 14353 21001
rect 13960 20967 14353 20968
rect 13960 20933 14289 20967
rect 14323 20933 14353 20967
rect 13960 20930 14353 20933
rect 13960 20896 14114 20930
rect 14148 20899 14353 20930
rect 14148 20896 14289 20899
rect 13960 20865 14289 20896
rect 14323 20865 14353 20899
rect 13960 20858 14353 20865
rect 13960 20824 14114 20858
rect 14148 20831 14353 20858
rect 14148 20824 14289 20831
rect 13960 20797 14289 20824
rect 14323 20797 14353 20831
rect 13960 20786 14353 20797
rect 13960 20752 14114 20786
rect 14148 20763 14353 20786
rect 14148 20752 14289 20763
rect 13960 20729 14289 20752
rect 14323 20729 14353 20763
rect 13960 20714 14353 20729
rect 13960 20680 14114 20714
rect 14148 20695 14353 20714
rect 14148 20680 14289 20695
rect 13960 20661 14289 20680
rect 14323 20661 14353 20695
rect 13960 20642 14353 20661
rect 13960 20608 14114 20642
rect 14148 20627 14353 20642
rect 14148 20608 14289 20627
rect 13960 20593 14289 20608
rect 14323 20593 14353 20627
rect 13960 20570 14353 20593
rect 13960 20536 14114 20570
rect 14148 20559 14353 20570
rect 14148 20536 14289 20559
rect 13960 20525 14289 20536
rect 14323 20525 14353 20559
rect 13960 20498 14353 20525
rect 13960 20464 14114 20498
rect 14148 20491 14353 20498
rect 14148 20464 14289 20491
rect 13960 20457 14289 20464
rect 14323 20457 14353 20491
rect 13960 20426 14353 20457
rect 13960 20392 14114 20426
rect 14148 20423 14353 20426
rect 14148 20392 14289 20423
rect 13960 20389 14289 20392
rect 14323 20389 14353 20423
rect 13960 20355 14353 20389
rect 13960 20354 14289 20355
rect 13960 20320 14114 20354
rect 14148 20321 14289 20354
rect 14323 20321 14353 20355
rect 14148 20320 14353 20321
rect 13960 20287 14353 20320
rect 13960 20282 14289 20287
rect 13960 20248 14114 20282
rect 14148 20253 14289 20282
rect 14323 20253 14353 20287
rect 14148 20248 14353 20253
rect 13960 20219 14353 20248
rect 13960 20210 14289 20219
rect 13960 20176 14114 20210
rect 14148 20185 14289 20210
rect 14323 20185 14353 20219
rect 14148 20176 14353 20185
rect 13960 20151 14353 20176
rect 13960 20138 14289 20151
rect 13960 20104 14114 20138
rect 14148 20117 14289 20138
rect 14323 20117 14353 20151
rect 14148 20104 14353 20117
rect 13960 20083 14353 20104
rect 13960 20066 14289 20083
rect 13960 20032 14114 20066
rect 14148 20049 14289 20066
rect 14323 20049 14353 20083
rect 14148 20032 14353 20049
rect 13960 20015 14353 20032
rect 13960 19994 14289 20015
rect 13960 19960 14114 19994
rect 14148 19981 14289 19994
rect 14323 19981 14353 20015
rect 14148 19960 14353 19981
rect 13960 19947 14353 19960
rect 13960 19922 14289 19947
rect 13960 19888 14114 19922
rect 14148 19913 14289 19922
rect 14323 19913 14353 19947
rect 14148 19888 14353 19913
rect 13960 19879 14353 19888
rect 13960 19850 14289 19879
rect 13960 19816 14114 19850
rect 14148 19845 14289 19850
rect 14323 19845 14353 19879
rect 14148 19816 14353 19845
rect 13960 19811 14353 19816
rect 13960 19778 14289 19811
rect 13960 19744 14114 19778
rect 14148 19777 14289 19778
rect 14323 19777 14353 19811
rect 14148 19744 14353 19777
rect 13960 19743 14353 19744
rect 13960 19709 14289 19743
rect 14323 19709 14353 19743
rect 13960 19706 14353 19709
rect 13960 19672 14114 19706
rect 14148 19675 14353 19706
rect 14148 19672 14289 19675
rect 13960 19641 14289 19672
rect 14323 19641 14353 19675
rect 13960 19634 14353 19641
rect 13960 19600 14114 19634
rect 14148 19607 14353 19634
rect 14148 19600 14289 19607
rect 13960 19573 14289 19600
rect 14323 19573 14353 19607
rect 13960 19562 14353 19573
rect 13960 19528 14114 19562
rect 14148 19539 14353 19562
rect 14148 19528 14289 19539
rect 13960 19505 14289 19528
rect 14323 19505 14353 19539
rect 13960 19490 14353 19505
rect 13960 19456 14114 19490
rect 14148 19471 14353 19490
rect 14148 19456 14289 19471
rect 13960 19437 14289 19456
rect 14323 19437 14353 19471
rect 13960 19418 14353 19437
rect 13960 19384 14114 19418
rect 14148 19403 14353 19418
rect 14148 19384 14289 19403
rect 13960 19369 14289 19384
rect 14323 19369 14353 19403
rect 13960 19346 14353 19369
rect 13960 19312 14114 19346
rect 14148 19335 14353 19346
rect 14148 19312 14289 19335
rect 13960 19301 14289 19312
rect 14323 19301 14353 19335
rect 13960 19274 14353 19301
rect 13960 19240 14114 19274
rect 14148 19267 14353 19274
rect 14148 19240 14289 19267
rect 13960 19233 14289 19240
rect 14323 19233 14353 19267
rect 13960 19202 14353 19233
rect 13960 19168 14114 19202
rect 14148 19199 14353 19202
rect 14148 19168 14289 19199
rect 13960 19165 14289 19168
rect 14323 19165 14353 19199
rect 13960 19131 14353 19165
rect 13960 19130 14289 19131
rect 13960 19096 14114 19130
rect 14148 19097 14289 19130
rect 14323 19097 14353 19131
rect 14148 19096 14353 19097
rect 13960 19063 14353 19096
rect 13960 19058 14289 19063
rect 13960 19024 14114 19058
rect 14148 19029 14289 19058
rect 14323 19029 14353 19063
rect 14148 19024 14353 19029
rect 13960 18995 14353 19024
rect 13960 18986 14289 18995
rect 13960 18952 14114 18986
rect 14148 18961 14289 18986
rect 14323 18961 14353 18995
rect 14148 18952 14353 18961
rect 13960 18927 14353 18952
rect 13960 18914 14289 18927
rect 13960 18880 14114 18914
rect 14148 18893 14289 18914
rect 14323 18893 14353 18927
rect 14148 18880 14353 18893
rect 13960 18859 14353 18880
rect 13960 18842 14289 18859
rect 13960 18808 14114 18842
rect 14148 18825 14289 18842
rect 14323 18825 14353 18859
rect 14148 18808 14353 18825
rect 13960 18791 14353 18808
rect 13960 18770 14289 18791
rect 13960 18736 14114 18770
rect 14148 18757 14289 18770
rect 14323 18757 14353 18791
rect 14148 18736 14353 18757
rect 13960 18723 14353 18736
rect 13960 18698 14289 18723
rect 13960 18664 14114 18698
rect 14148 18689 14289 18698
rect 14323 18689 14353 18723
rect 14148 18664 14353 18689
rect 13960 18655 14353 18664
rect 13960 18626 14289 18655
rect 13960 18592 14114 18626
rect 14148 18621 14289 18626
rect 14323 18621 14353 18655
rect 14148 18592 14353 18621
rect 13960 18587 14353 18592
rect 13960 18554 14289 18587
rect 13960 18520 14114 18554
rect 14148 18553 14289 18554
rect 14323 18553 14353 18587
rect 14148 18520 14353 18553
rect 13960 18519 14353 18520
rect 13960 18485 14289 18519
rect 14323 18485 14353 18519
rect 13960 18482 14353 18485
rect 13960 18448 14114 18482
rect 14148 18451 14353 18482
rect 14148 18448 14289 18451
rect 13960 18417 14289 18448
rect 14323 18417 14353 18451
rect 13960 18410 14353 18417
rect 13960 18376 14114 18410
rect 14148 18383 14353 18410
rect 14148 18376 14289 18383
rect 13960 18349 14289 18376
rect 14323 18349 14353 18383
rect 13960 18338 14353 18349
rect 13960 18304 14114 18338
rect 14148 18315 14353 18338
rect 14148 18304 14289 18315
rect 13960 18281 14289 18304
rect 14323 18281 14353 18315
rect 13960 18266 14353 18281
rect 13960 18232 14114 18266
rect 14148 18247 14353 18266
rect 14148 18232 14289 18247
rect 13960 18213 14289 18232
rect 14323 18213 14353 18247
rect 13960 18194 14353 18213
rect 13960 18160 14114 18194
rect 14148 18179 14353 18194
rect 14148 18160 14289 18179
rect 13960 18145 14289 18160
rect 14323 18145 14353 18179
rect 13960 18122 14353 18145
rect 13960 18088 14114 18122
rect 14148 18111 14353 18122
rect 14148 18088 14289 18111
rect 13960 18077 14289 18088
rect 14323 18077 14353 18111
rect 13960 18050 14353 18077
rect 13960 18016 14114 18050
rect 14148 18043 14353 18050
rect 14148 18016 14289 18043
rect 13960 18009 14289 18016
rect 14323 18009 14353 18043
rect 13960 17978 14353 18009
rect 13960 17944 14114 17978
rect 14148 17975 14353 17978
rect 14148 17944 14289 17975
rect 13960 17941 14289 17944
rect 14323 17941 14353 17975
rect 13960 17907 14353 17941
rect 13960 17906 14289 17907
rect 13960 17872 14114 17906
rect 14148 17873 14289 17906
rect 14323 17873 14353 17907
rect 14148 17872 14353 17873
rect 13960 17839 14353 17872
rect 13960 17834 14289 17839
rect 13960 17800 14114 17834
rect 14148 17805 14289 17834
rect 14323 17805 14353 17839
rect 14148 17800 14353 17805
rect 13960 17771 14353 17800
rect 13960 17762 14289 17771
rect 13960 17728 14114 17762
rect 14148 17737 14289 17762
rect 14323 17737 14353 17771
rect 14148 17728 14353 17737
rect 13960 17703 14353 17728
rect 13960 17690 14289 17703
rect 13960 17656 14114 17690
rect 14148 17669 14289 17690
rect 14323 17669 14353 17703
rect 14148 17656 14353 17669
rect 13960 17635 14353 17656
rect 13960 17618 14289 17635
rect 13960 17584 14114 17618
rect 14148 17601 14289 17618
rect 14323 17601 14353 17635
rect 14148 17584 14353 17601
rect 13960 17567 14353 17584
rect 13960 17546 14289 17567
rect 13960 17512 14114 17546
rect 14148 17533 14289 17546
rect 14323 17533 14353 17567
rect 14148 17512 14353 17533
rect 13960 17499 14353 17512
rect 13960 17474 14289 17499
rect 13960 17440 14114 17474
rect 14148 17465 14289 17474
rect 14323 17465 14353 17499
rect 14148 17440 14353 17465
rect 13960 17431 14353 17440
rect 13960 17402 14289 17431
rect 13960 17368 14114 17402
rect 14148 17397 14289 17402
rect 14323 17397 14353 17431
rect 14148 17368 14353 17397
rect 13960 17363 14353 17368
rect 13960 17330 14289 17363
rect 13960 17296 14114 17330
rect 14148 17329 14289 17330
rect 14323 17329 14353 17363
rect 14148 17296 14353 17329
rect 13960 17295 14353 17296
rect 13960 17261 14289 17295
rect 14323 17261 14353 17295
rect 13960 17258 14353 17261
rect 13960 17224 14114 17258
rect 14148 17227 14353 17258
rect 14148 17224 14289 17227
rect 13960 17193 14289 17224
rect 14323 17193 14353 17227
rect 13960 17186 14353 17193
rect 13960 17152 14114 17186
rect 14148 17159 14353 17186
rect 14148 17152 14289 17159
rect 13960 17125 14289 17152
rect 14323 17125 14353 17159
rect 13960 17114 14353 17125
rect 13960 17080 14114 17114
rect 14148 17091 14353 17114
rect 14148 17080 14289 17091
rect 13960 17057 14289 17080
rect 14323 17057 14353 17091
rect 13960 17042 14353 17057
rect 13960 17008 14114 17042
rect 14148 17023 14353 17042
rect 14148 17008 14289 17023
rect 13960 16989 14289 17008
rect 14323 16989 14353 17023
rect 13960 16970 14353 16989
rect 13960 16936 14114 16970
rect 14148 16955 14353 16970
rect 14148 16936 14289 16955
rect 13960 16921 14289 16936
rect 14323 16921 14353 16955
rect 13960 16898 14353 16921
rect 13960 16864 14114 16898
rect 14148 16887 14353 16898
rect 14148 16864 14289 16887
rect 13960 16853 14289 16864
rect 14323 16853 14353 16887
rect 13960 16826 14353 16853
rect 13960 16792 14114 16826
rect 14148 16819 14353 16826
rect 14148 16792 14289 16819
rect 13960 16785 14289 16792
rect 14323 16785 14353 16819
rect 13960 16754 14353 16785
rect 13960 16720 14114 16754
rect 14148 16751 14353 16754
rect 14148 16720 14289 16751
rect 13960 16717 14289 16720
rect 14323 16717 14353 16751
rect 13960 16683 14353 16717
rect 13960 16682 14289 16683
rect 13960 16648 14114 16682
rect 14148 16649 14289 16682
rect 14323 16649 14353 16683
rect 14148 16648 14353 16649
rect 13960 16615 14353 16648
rect 13960 16610 14289 16615
rect 13960 16576 14114 16610
rect 14148 16581 14289 16610
rect 14323 16581 14353 16615
rect 14148 16576 14353 16581
rect 13960 16547 14353 16576
rect 13960 16538 14289 16547
rect 13960 16504 14114 16538
rect 14148 16513 14289 16538
rect 14323 16513 14353 16547
rect 14148 16504 14353 16513
rect 13960 16479 14353 16504
rect 13960 16466 14289 16479
rect 13960 16432 14114 16466
rect 14148 16445 14289 16466
rect 14323 16445 14353 16479
rect 14148 16432 14353 16445
rect 13960 16411 14353 16432
rect 13960 16394 14289 16411
rect 13960 16360 14114 16394
rect 14148 16377 14289 16394
rect 14323 16377 14353 16411
rect 14148 16360 14353 16377
rect 13960 16343 14353 16360
rect 13960 16322 14289 16343
rect 13960 16288 14114 16322
rect 14148 16309 14289 16322
rect 14323 16309 14353 16343
rect 14148 16288 14353 16309
rect 13960 16275 14353 16288
rect 13960 16250 14289 16275
rect 13960 16216 14114 16250
rect 14148 16241 14289 16250
rect 14323 16241 14353 16275
rect 14148 16216 14353 16241
rect 13960 16207 14353 16216
rect 13960 16178 14289 16207
rect 13960 16144 14114 16178
rect 14148 16173 14289 16178
rect 14323 16173 14353 16207
rect 14148 16144 14353 16173
rect 13960 16139 14353 16144
rect 13960 16106 14289 16139
rect 13960 16072 14114 16106
rect 14148 16105 14289 16106
rect 14323 16105 14353 16139
rect 14148 16072 14353 16105
rect 13960 16071 14353 16072
rect 13960 16037 14289 16071
rect 14323 16037 14353 16071
rect 13960 16034 14353 16037
rect 13960 16000 14114 16034
rect 14148 16003 14353 16034
rect 14148 16000 14289 16003
rect 13960 15969 14289 16000
rect 14323 15969 14353 16003
rect 13960 15962 14353 15969
rect 13960 15928 14114 15962
rect 14148 15935 14353 15962
rect 14148 15928 14289 15935
rect 13960 15901 14289 15928
rect 14323 15901 14353 15935
rect 13960 15890 14353 15901
rect 13960 15856 14114 15890
rect 14148 15867 14353 15890
rect 14148 15856 14289 15867
rect 13960 15833 14289 15856
rect 14323 15833 14353 15867
rect 13960 15818 14353 15833
rect 13960 15784 14114 15818
rect 14148 15799 14353 15818
rect 14148 15784 14289 15799
rect 13960 15765 14289 15784
rect 14323 15765 14353 15799
rect 13960 15746 14353 15765
rect 13960 15712 14114 15746
rect 14148 15731 14353 15746
rect 14148 15712 14289 15731
rect 13960 15697 14289 15712
rect 14323 15697 14353 15731
rect 13960 15674 14353 15697
rect 13960 15640 14114 15674
rect 14148 15663 14353 15674
rect 14148 15640 14289 15663
rect 13960 15629 14289 15640
rect 14323 15629 14353 15663
rect 13960 15602 14353 15629
rect 13960 15568 14114 15602
rect 14148 15595 14353 15602
rect 14148 15568 14289 15595
rect 13960 15561 14289 15568
rect 14323 15561 14353 15595
rect 13960 15530 14353 15561
rect 13960 15496 14114 15530
rect 14148 15527 14353 15530
rect 14148 15496 14289 15527
rect 13960 15493 14289 15496
rect 14323 15493 14353 15527
rect 13960 15459 14353 15493
rect 13960 15458 14289 15459
rect 13960 15424 14114 15458
rect 14148 15425 14289 15458
rect 14323 15425 14353 15459
rect 14148 15424 14353 15425
rect 13960 15391 14353 15424
rect 13960 15386 14289 15391
rect 13960 15352 14114 15386
rect 14148 15357 14289 15386
rect 14323 15357 14353 15391
rect 14148 15352 14353 15357
rect 13960 15323 14353 15352
rect 13960 15314 14289 15323
rect 13960 15280 14114 15314
rect 14148 15289 14289 15314
rect 14323 15289 14353 15323
rect 14148 15280 14353 15289
rect 13960 15255 14353 15280
rect 13960 15242 14289 15255
rect 595 15153 624 15187
rect 658 15177 1018 15187
rect 658 15153 799 15177
rect 595 15143 799 15153
rect 833 15143 1018 15177
rect 595 15119 1018 15143
rect 595 15085 624 15119
rect 658 15105 1018 15119
rect 658 15085 799 15105
rect 595 15071 799 15085
rect 833 15101 1018 15105
rect 13960 15208 14114 15242
rect 14148 15221 14289 15242
rect 14323 15221 14353 15255
rect 14148 15208 14353 15221
rect 13960 15187 14353 15208
rect 13960 15170 14289 15187
rect 13960 15136 14114 15170
rect 14148 15153 14289 15170
rect 14323 15153 14353 15187
rect 14148 15136 14353 15153
rect 13960 15119 14353 15136
rect 13960 15101 14289 15119
rect 833 15098 14289 15101
rect 833 15071 14114 15098
rect 595 15064 14114 15071
rect 14148 15085 14289 15098
rect 14323 15085 14353 15119
rect 14148 15064 14353 15085
rect 595 15051 14353 15064
rect 595 15017 624 15051
rect 658 15017 14289 15051
rect 14323 15017 14353 15051
rect 595 14983 14353 15017
rect 595 14949 624 14983
rect 658 14955 14289 14983
rect 658 14949 883 14955
rect 595 14921 883 14949
rect 917 14921 955 14955
rect 989 14921 1027 14955
rect 1061 14921 1099 14955
rect 1133 14921 1171 14955
rect 1205 14921 1243 14955
rect 1277 14921 1315 14955
rect 1349 14921 1387 14955
rect 1421 14921 1459 14955
rect 1493 14921 1531 14955
rect 1565 14921 1603 14955
rect 1637 14921 1675 14955
rect 1709 14921 1747 14955
rect 1781 14921 1819 14955
rect 1853 14921 1891 14955
rect 1925 14921 1963 14955
rect 1997 14921 2035 14955
rect 2069 14921 2107 14955
rect 2141 14921 2179 14955
rect 2213 14921 2251 14955
rect 2285 14921 2323 14955
rect 2357 14921 2395 14955
rect 2429 14921 2467 14955
rect 2501 14921 2539 14955
rect 2573 14921 2611 14955
rect 2645 14921 2683 14955
rect 2717 14921 2755 14955
rect 2789 14921 2827 14955
rect 2861 14921 2899 14955
rect 2933 14921 2971 14955
rect 3005 14921 3043 14955
rect 3077 14921 3115 14955
rect 3149 14921 3187 14955
rect 3221 14921 3259 14955
rect 3293 14921 3331 14955
rect 3365 14921 3403 14955
rect 3437 14921 3475 14955
rect 3509 14921 3547 14955
rect 3581 14921 3619 14955
rect 3653 14921 3691 14955
rect 3725 14921 3763 14955
rect 3797 14921 3835 14955
rect 3869 14921 3907 14955
rect 3941 14921 3979 14955
rect 4013 14921 4051 14955
rect 4085 14921 4123 14955
rect 4157 14921 4195 14955
rect 4229 14921 4267 14955
rect 4301 14921 4339 14955
rect 4373 14921 4411 14955
rect 4445 14921 4483 14955
rect 4517 14921 4555 14955
rect 4589 14921 4627 14955
rect 4661 14921 4699 14955
rect 4733 14921 4771 14955
rect 4805 14921 4843 14955
rect 4877 14921 4915 14955
rect 4949 14921 4987 14955
rect 5021 14921 5059 14955
rect 5093 14921 5131 14955
rect 5165 14921 5203 14955
rect 5237 14921 5275 14955
rect 5309 14921 5347 14955
rect 5381 14921 5419 14955
rect 5453 14921 5491 14955
rect 5525 14921 5563 14955
rect 5597 14921 5635 14955
rect 5669 14921 5707 14955
rect 5741 14921 5779 14955
rect 5813 14921 5851 14955
rect 5885 14921 5923 14955
rect 5957 14921 5995 14955
rect 6029 14921 6067 14955
rect 6101 14921 6139 14955
rect 6173 14921 6211 14955
rect 6245 14921 6283 14955
rect 6317 14921 6355 14955
rect 6389 14921 6427 14955
rect 6461 14921 6499 14955
rect 6533 14921 6571 14955
rect 6605 14921 6643 14955
rect 6677 14921 6715 14955
rect 6749 14921 6787 14955
rect 6821 14921 6859 14955
rect 6893 14921 6931 14955
rect 6965 14921 7003 14955
rect 7037 14921 7075 14955
rect 7109 14921 7147 14955
rect 7181 14921 7219 14955
rect 7253 14921 7291 14955
rect 7325 14921 7363 14955
rect 7397 14921 7435 14955
rect 7469 14921 7507 14955
rect 7541 14921 7579 14955
rect 7613 14921 7651 14955
rect 7685 14921 7723 14955
rect 7757 14921 7795 14955
rect 7829 14921 7867 14955
rect 7901 14921 7939 14955
rect 7973 14921 8011 14955
rect 8045 14921 8083 14955
rect 8117 14921 8155 14955
rect 8189 14921 8227 14955
rect 8261 14921 8299 14955
rect 8333 14921 8371 14955
rect 8405 14921 8443 14955
rect 8477 14921 8515 14955
rect 8549 14921 8587 14955
rect 8621 14921 8659 14955
rect 8693 14921 8731 14955
rect 8765 14921 8803 14955
rect 8837 14921 8875 14955
rect 8909 14921 8947 14955
rect 8981 14921 9019 14955
rect 9053 14921 9091 14955
rect 9125 14921 9163 14955
rect 9197 14921 9235 14955
rect 9269 14921 9307 14955
rect 9341 14921 9379 14955
rect 9413 14921 9451 14955
rect 9485 14921 9523 14955
rect 9557 14921 9595 14955
rect 9629 14921 9667 14955
rect 9701 14921 9739 14955
rect 9773 14921 9811 14955
rect 9845 14921 9883 14955
rect 9917 14921 9955 14955
rect 9989 14921 10027 14955
rect 10061 14921 10099 14955
rect 10133 14921 10171 14955
rect 10205 14921 10243 14955
rect 10277 14921 10315 14955
rect 10349 14921 10387 14955
rect 10421 14921 10459 14955
rect 10493 14921 10531 14955
rect 10565 14921 10603 14955
rect 10637 14921 10675 14955
rect 10709 14921 10747 14955
rect 10781 14921 10819 14955
rect 10853 14921 10891 14955
rect 10925 14921 10963 14955
rect 10997 14921 11035 14955
rect 11069 14921 11107 14955
rect 11141 14921 11179 14955
rect 11213 14921 11251 14955
rect 11285 14921 11323 14955
rect 11357 14921 11395 14955
rect 11429 14921 11467 14955
rect 11501 14921 11539 14955
rect 11573 14921 11611 14955
rect 11645 14921 11683 14955
rect 11717 14921 11755 14955
rect 11789 14921 11827 14955
rect 11861 14921 11899 14955
rect 11933 14921 11971 14955
rect 12005 14921 12043 14955
rect 12077 14921 12115 14955
rect 12149 14921 12187 14955
rect 12221 14921 12259 14955
rect 12293 14921 12331 14955
rect 12365 14921 12403 14955
rect 12437 14921 12475 14955
rect 12509 14921 12547 14955
rect 12581 14921 12619 14955
rect 12653 14921 12691 14955
rect 12725 14921 12763 14955
rect 12797 14921 12835 14955
rect 12869 14921 12907 14955
rect 12941 14921 12979 14955
rect 13013 14921 13051 14955
rect 13085 14921 13123 14955
rect 13157 14921 13195 14955
rect 13229 14921 13267 14955
rect 13301 14921 13339 14955
rect 13373 14921 13411 14955
rect 13445 14921 13483 14955
rect 13517 14921 13555 14955
rect 13589 14921 13627 14955
rect 13661 14921 13699 14955
rect 13733 14921 13771 14955
rect 13805 14921 13843 14955
rect 13877 14921 13915 14955
rect 13949 14921 13987 14955
rect 14021 14949 14289 14955
rect 14323 14949 14353 14983
rect 14021 14921 14353 14949
rect 595 14915 14353 14921
rect 595 14881 624 14915
rect 658 14881 14289 14915
rect 14323 14881 14353 14915
rect 595 14788 14353 14881
rect 595 14754 758 14788
rect 792 14754 826 14788
rect 860 14787 894 14788
rect 928 14787 962 14788
rect 996 14787 1030 14788
rect 1064 14787 1098 14788
rect 1132 14787 1166 14788
rect 860 14754 875 14787
rect 928 14754 947 14787
rect 996 14754 1019 14787
rect 1064 14754 1091 14787
rect 1132 14754 1163 14787
rect 1200 14754 1234 14788
rect 1268 14787 1302 14788
rect 1336 14787 1370 14788
rect 1404 14787 1438 14788
rect 1472 14787 1506 14788
rect 1540 14787 1574 14788
rect 1608 14787 1642 14788
rect 1676 14787 1710 14788
rect 1744 14787 1778 14788
rect 1812 14787 1846 14788
rect 1269 14754 1302 14787
rect 1341 14754 1370 14787
rect 1413 14754 1438 14787
rect 1485 14754 1506 14787
rect 1557 14754 1574 14787
rect 1629 14754 1642 14787
rect 1701 14754 1710 14787
rect 1773 14754 1778 14787
rect 1845 14754 1846 14787
rect 1880 14787 1914 14788
rect 1948 14787 1982 14788
rect 2016 14787 2050 14788
rect 1880 14754 1883 14787
rect 1948 14754 1955 14787
rect 2016 14754 2027 14787
rect 2084 14754 2118 14788
rect 2152 14754 2186 14788
rect 2220 14754 2254 14788
rect 2288 14754 2322 14788
rect 2356 14754 2390 14788
rect 2424 14754 2458 14788
rect 2492 14754 2526 14788
rect 2560 14754 2594 14788
rect 2628 14754 2662 14788
rect 2696 14754 2730 14788
rect 2764 14754 2798 14788
rect 2832 14754 2866 14788
rect 2900 14754 2934 14788
rect 2968 14754 3002 14788
rect 3036 14754 3070 14788
rect 3104 14754 3138 14788
rect 3172 14754 3206 14788
rect 3240 14754 3274 14788
rect 3308 14754 3342 14788
rect 3376 14754 3410 14788
rect 3444 14754 3478 14788
rect 3512 14754 3546 14788
rect 3580 14754 3614 14788
rect 3648 14754 3682 14788
rect 3716 14754 3750 14788
rect 3784 14754 3818 14788
rect 3852 14754 3886 14788
rect 3920 14754 3954 14788
rect 3988 14754 4022 14788
rect 4056 14754 4090 14788
rect 4124 14754 4158 14788
rect 4192 14754 4226 14788
rect 4260 14754 4294 14788
rect 4328 14754 4362 14788
rect 4396 14754 4430 14788
rect 4464 14754 4498 14788
rect 4532 14754 4566 14788
rect 4600 14754 4634 14788
rect 4668 14754 4702 14788
rect 4736 14754 4770 14788
rect 4804 14754 4838 14788
rect 4872 14754 4906 14788
rect 4940 14754 4974 14788
rect 5008 14754 5042 14788
rect 5076 14754 5110 14788
rect 5144 14754 5178 14788
rect 5212 14754 5246 14788
rect 5280 14754 5314 14788
rect 5348 14754 5382 14788
rect 5416 14754 5450 14788
rect 5484 14754 5518 14788
rect 5552 14754 5586 14788
rect 5620 14754 5654 14788
rect 5688 14754 5722 14788
rect 5756 14754 5790 14788
rect 5824 14754 5858 14788
rect 5892 14754 5926 14788
rect 5960 14754 5994 14788
rect 6028 14754 6062 14788
rect 6096 14754 6130 14788
rect 6164 14754 6198 14788
rect 6232 14754 6266 14788
rect 6300 14754 6334 14788
rect 6368 14754 6402 14788
rect 6436 14754 6470 14788
rect 6504 14754 6538 14788
rect 6572 14754 6606 14788
rect 6640 14754 6674 14788
rect 6708 14754 6742 14788
rect 6776 14754 6810 14788
rect 6844 14754 6878 14788
rect 6912 14754 6946 14788
rect 6980 14754 7014 14788
rect 7048 14754 7082 14788
rect 7116 14754 7150 14788
rect 7184 14754 7218 14788
rect 7252 14754 7286 14788
rect 7320 14754 7354 14788
rect 7388 14754 7422 14788
rect 7456 14754 7490 14788
rect 7524 14754 7558 14788
rect 7592 14754 7626 14788
rect 7660 14754 7694 14788
rect 7728 14754 7762 14788
rect 7796 14754 7830 14788
rect 7864 14754 7898 14788
rect 7932 14754 7966 14788
rect 8000 14754 8034 14788
rect 8068 14754 8102 14788
rect 8136 14754 8170 14788
rect 8204 14754 8238 14788
rect 8272 14754 8306 14788
rect 8340 14754 8374 14788
rect 8408 14754 8442 14788
rect 8476 14754 8510 14788
rect 8544 14754 8578 14788
rect 8612 14754 8646 14788
rect 8680 14754 8714 14788
rect 8748 14754 8782 14788
rect 8816 14754 8850 14788
rect 8884 14754 8918 14788
rect 8952 14754 8986 14788
rect 9020 14754 9054 14788
rect 9088 14754 9122 14788
rect 9156 14754 9190 14788
rect 9224 14754 9258 14788
rect 9292 14754 9326 14788
rect 9360 14754 9394 14788
rect 9428 14754 9462 14788
rect 9496 14754 9530 14788
rect 9564 14754 9598 14788
rect 9632 14754 9666 14788
rect 9700 14754 9734 14788
rect 9768 14754 9802 14788
rect 9836 14754 9870 14788
rect 9904 14754 9938 14788
rect 9972 14754 10006 14788
rect 10040 14754 10074 14788
rect 10108 14754 10142 14788
rect 10176 14754 10210 14788
rect 10244 14754 10278 14788
rect 10312 14754 10346 14788
rect 10380 14754 10414 14788
rect 10448 14754 10482 14788
rect 10516 14754 10550 14788
rect 10584 14754 10618 14788
rect 10652 14754 10686 14788
rect 10720 14754 10754 14788
rect 10788 14754 10822 14788
rect 10856 14754 10890 14788
rect 10924 14754 10958 14788
rect 10992 14754 11026 14788
rect 11060 14754 11094 14788
rect 11128 14754 11162 14788
rect 11196 14754 11230 14788
rect 11264 14754 11298 14788
rect 11332 14754 11366 14788
rect 11400 14754 11434 14788
rect 11468 14754 11502 14788
rect 11536 14754 11570 14788
rect 11604 14754 11638 14788
rect 11672 14754 11706 14788
rect 11740 14754 11774 14788
rect 11808 14754 11842 14788
rect 11876 14754 11910 14788
rect 11944 14754 11978 14788
rect 12012 14754 12046 14788
rect 12080 14754 12114 14788
rect 12148 14754 12182 14788
rect 12216 14754 12250 14788
rect 12284 14754 12318 14788
rect 12352 14754 12386 14788
rect 12420 14754 12454 14788
rect 12488 14754 12522 14788
rect 12556 14754 12590 14788
rect 12624 14754 12658 14788
rect 12692 14754 12726 14788
rect 12760 14754 12794 14788
rect 12828 14754 12862 14788
rect 12896 14787 12930 14788
rect 12964 14787 12998 14788
rect 13032 14787 13066 14788
rect 13100 14787 13134 14788
rect 13168 14787 13202 14788
rect 13236 14787 13270 14788
rect 12909 14754 12930 14787
rect 12981 14754 12998 14787
rect 13053 14754 13066 14787
rect 13125 14754 13134 14787
rect 13197 14754 13202 14787
rect 13269 14754 13270 14787
rect 13304 14787 13338 14788
rect 13372 14787 13406 14788
rect 13440 14787 13474 14788
rect 13508 14787 13542 14788
rect 13576 14787 13610 14788
rect 13644 14787 13678 14788
rect 13712 14787 13746 14788
rect 13780 14787 13814 14788
rect 13304 14754 13307 14787
rect 13372 14754 13379 14787
rect 13440 14754 13451 14787
rect 13508 14754 13523 14787
rect 13576 14754 13595 14787
rect 13644 14754 13667 14787
rect 13712 14754 13739 14787
rect 13780 14754 13811 14787
rect 13848 14754 13882 14788
rect 13916 14787 13950 14788
rect 13984 14787 14018 14788
rect 14052 14787 14086 14788
rect 13917 14754 13950 14787
rect 13989 14754 14018 14787
rect 14061 14754 14086 14787
rect 14120 14754 14154 14788
rect 14188 14754 14353 14788
rect 595 14753 875 14754
rect 909 14753 947 14754
rect 981 14753 1019 14754
rect 1053 14753 1091 14754
rect 1125 14753 1163 14754
rect 1197 14753 1235 14754
rect 1269 14753 1307 14754
rect 1341 14753 1379 14754
rect 1413 14753 1451 14754
rect 1485 14753 1523 14754
rect 1557 14753 1595 14754
rect 1629 14753 1667 14754
rect 1701 14753 1739 14754
rect 1773 14753 1811 14754
rect 1845 14753 1883 14754
rect 1917 14753 1955 14754
rect 1989 14753 2027 14754
rect 2061 14753 12875 14754
rect 12909 14753 12947 14754
rect 12981 14753 13019 14754
rect 13053 14753 13091 14754
rect 13125 14753 13163 14754
rect 13197 14753 13235 14754
rect 13269 14753 13307 14754
rect 13341 14753 13379 14754
rect 13413 14753 13451 14754
rect 13485 14753 13523 14754
rect 13557 14753 13595 14754
rect 13629 14753 13667 14754
rect 13701 14753 13739 14754
rect 13773 14753 13811 14754
rect 13845 14753 13883 14754
rect 13917 14753 13955 14754
rect 13989 14753 14027 14754
rect 14061 14753 14353 14754
rect 595 14724 14353 14753
rect 14531 36205 14599 36239
rect 14633 36219 14716 36239
rect 14531 36185 14606 36205
rect 14640 36185 14716 36219
rect 14531 36171 14716 36185
rect 14531 36137 14599 36171
rect 14633 36147 14716 36171
rect 14531 36113 14606 36137
rect 14640 36113 14716 36147
rect 14531 36103 14716 36113
rect 14531 36069 14599 36103
rect 14633 36075 14716 36103
rect 14531 36041 14606 36069
rect 14640 36041 14716 36075
rect 14531 36035 14716 36041
rect 14531 36001 14599 36035
rect 14633 36003 14716 36035
rect 14531 35969 14606 36001
rect 14640 35969 14716 36003
rect 14531 35967 14716 35969
rect 14531 35933 14599 35967
rect 14633 35933 14716 35967
rect 14531 35931 14716 35933
rect 14531 35899 14606 35931
rect 14531 35865 14599 35899
rect 14640 35897 14716 35931
rect 14633 35865 14716 35897
rect 14531 35859 14716 35865
rect 14531 35831 14606 35859
rect 14531 35797 14599 35831
rect 14640 35825 14716 35859
rect 14633 35797 14716 35825
rect 14531 35787 14716 35797
rect 14531 35763 14606 35787
rect 14531 35729 14599 35763
rect 14640 35753 14716 35787
rect 14633 35729 14716 35753
rect 14531 35715 14716 35729
rect 14531 35695 14606 35715
rect 14531 35661 14599 35695
rect 14640 35681 14716 35715
rect 14633 35661 14716 35681
rect 14531 35643 14716 35661
rect 14531 35627 14606 35643
rect 14531 35593 14599 35627
rect 14640 35609 14716 35643
rect 14633 35593 14716 35609
rect 14531 35571 14716 35593
rect 14531 35559 14606 35571
rect 14531 35525 14599 35559
rect 14640 35537 14716 35571
rect 14633 35525 14716 35537
rect 14531 35499 14716 35525
rect 14531 35491 14606 35499
rect 14531 35457 14599 35491
rect 14640 35465 14716 35499
rect 14633 35457 14716 35465
rect 14531 35427 14716 35457
rect 14531 35423 14606 35427
rect 14531 35389 14599 35423
rect 14640 35393 14716 35427
rect 14633 35389 14716 35393
rect 14531 35355 14716 35389
rect 14531 35321 14599 35355
rect 14640 35321 14716 35355
rect 14531 35287 14716 35321
rect 14531 35253 14599 35287
rect 14633 35283 14716 35287
rect 14531 35249 14606 35253
rect 14640 35249 14716 35283
rect 14531 35219 14716 35249
rect 14531 35185 14599 35219
rect 14633 35211 14716 35219
rect 14531 35177 14606 35185
rect 14640 35177 14716 35211
rect 14531 35151 14716 35177
rect 14531 35117 14599 35151
rect 14633 35139 14716 35151
rect 14531 35105 14606 35117
rect 14640 35105 14716 35139
rect 14531 35083 14716 35105
rect 14531 35049 14599 35083
rect 14633 35067 14716 35083
rect 14531 35033 14606 35049
rect 14640 35033 14716 35067
rect 14531 35015 14716 35033
rect 14531 34981 14599 35015
rect 14633 34995 14716 35015
rect 14531 34961 14606 34981
rect 14640 34961 14716 34995
rect 14531 34947 14716 34961
rect 14531 34913 14599 34947
rect 14633 34923 14716 34947
rect 14531 34889 14606 34913
rect 14640 34889 14716 34923
rect 14531 34879 14716 34889
rect 14531 34845 14599 34879
rect 14633 34851 14716 34879
rect 14531 34817 14606 34845
rect 14640 34817 14716 34851
rect 14531 34811 14716 34817
rect 14531 34777 14599 34811
rect 14633 34779 14716 34811
rect 14531 34745 14606 34777
rect 14640 34745 14716 34779
rect 14531 34743 14716 34745
rect 14531 34709 14599 34743
rect 14633 34709 14716 34743
rect 14531 34707 14716 34709
rect 14531 34675 14606 34707
rect 14531 34641 14599 34675
rect 14640 34673 14716 34707
rect 14633 34641 14716 34673
rect 14531 34635 14716 34641
rect 14531 34607 14606 34635
rect 14531 34573 14599 34607
rect 14640 34601 14716 34635
rect 14633 34573 14716 34601
rect 14531 34563 14716 34573
rect 14531 34539 14606 34563
rect 14531 34505 14599 34539
rect 14640 34529 14716 34563
rect 14633 34505 14716 34529
rect 14531 34491 14716 34505
rect 14531 34471 14606 34491
rect 14531 34437 14599 34471
rect 14640 34457 14716 34491
rect 14633 34437 14716 34457
rect 14531 34419 14716 34437
rect 14531 34403 14606 34419
rect 14531 34369 14599 34403
rect 14640 34385 14716 34419
rect 14633 34369 14716 34385
rect 14531 34347 14716 34369
rect 14531 34335 14606 34347
rect 14531 34301 14599 34335
rect 14640 34313 14716 34347
rect 14633 34301 14716 34313
rect 14531 34275 14716 34301
rect 14531 34267 14606 34275
rect 14531 34233 14599 34267
rect 14640 34241 14716 34275
rect 14633 34233 14716 34241
rect 14531 34203 14716 34233
rect 14531 34199 14606 34203
rect 14531 34165 14599 34199
rect 14640 34169 14716 34203
rect 14633 34165 14716 34169
rect 14531 34131 14716 34165
rect 14531 34097 14599 34131
rect 14640 34097 14716 34131
rect 14531 34063 14716 34097
rect 14531 34029 14599 34063
rect 14633 34059 14716 34063
rect 14531 34025 14606 34029
rect 14640 34025 14716 34059
rect 14531 33995 14716 34025
rect 14531 33961 14599 33995
rect 14633 33987 14716 33995
rect 14531 33953 14606 33961
rect 14640 33953 14716 33987
rect 14531 33927 14716 33953
rect 14531 33893 14599 33927
rect 14633 33915 14716 33927
rect 14531 33881 14606 33893
rect 14640 33881 14716 33915
rect 14531 33859 14716 33881
rect 14531 33825 14599 33859
rect 14633 33843 14716 33859
rect 14531 33809 14606 33825
rect 14640 33809 14716 33843
rect 14531 33791 14716 33809
rect 14531 33757 14599 33791
rect 14633 33771 14716 33791
rect 14531 33737 14606 33757
rect 14640 33737 14716 33771
rect 14531 33723 14716 33737
rect 14531 33689 14599 33723
rect 14633 33699 14716 33723
rect 14531 33665 14606 33689
rect 14640 33665 14716 33699
rect 14531 33655 14716 33665
rect 14531 33621 14599 33655
rect 14633 33627 14716 33655
rect 14531 33593 14606 33621
rect 14640 33593 14716 33627
rect 14531 33587 14716 33593
rect 14531 33553 14599 33587
rect 14633 33555 14716 33587
rect 14531 33521 14606 33553
rect 14640 33521 14716 33555
rect 14531 33519 14716 33521
rect 14531 33485 14599 33519
rect 14633 33485 14716 33519
rect 14531 33483 14716 33485
rect 14531 33451 14606 33483
rect 14531 33417 14599 33451
rect 14640 33449 14716 33483
rect 14633 33417 14716 33449
rect 14531 33411 14716 33417
rect 14531 33383 14606 33411
rect 14531 33349 14599 33383
rect 14640 33377 14716 33411
rect 14633 33349 14716 33377
rect 14531 33339 14716 33349
rect 14531 33315 14606 33339
rect 14531 33281 14599 33315
rect 14640 33305 14716 33339
rect 14633 33281 14716 33305
rect 14531 33267 14716 33281
rect 14531 33247 14606 33267
rect 14531 33213 14599 33247
rect 14640 33233 14716 33267
rect 14633 33213 14716 33233
rect 14531 33195 14716 33213
rect 14531 33179 14606 33195
rect 14531 33145 14599 33179
rect 14640 33161 14716 33195
rect 14633 33145 14716 33161
rect 14531 33123 14716 33145
rect 14531 33111 14606 33123
rect 14531 33077 14599 33111
rect 14640 33089 14716 33123
rect 14633 33077 14716 33089
rect 14531 33051 14716 33077
rect 14531 33043 14606 33051
rect 14531 33009 14599 33043
rect 14640 33017 14716 33051
rect 14633 33009 14716 33017
rect 14531 32979 14716 33009
rect 14531 32975 14606 32979
rect 14531 32941 14599 32975
rect 14640 32945 14716 32979
rect 14633 32941 14716 32945
rect 14531 32907 14716 32941
rect 14531 32873 14599 32907
rect 14640 32873 14716 32907
rect 14531 32839 14716 32873
rect 14531 32805 14599 32839
rect 14633 32835 14716 32839
rect 14531 32801 14606 32805
rect 14640 32801 14716 32835
rect 14531 32771 14716 32801
rect 14531 32737 14599 32771
rect 14633 32763 14716 32771
rect 14531 32729 14606 32737
rect 14640 32729 14716 32763
rect 14531 32703 14716 32729
rect 14531 32669 14599 32703
rect 14633 32691 14716 32703
rect 14531 32657 14606 32669
rect 14640 32657 14716 32691
rect 14531 32635 14716 32657
rect 14531 32601 14599 32635
rect 14633 32619 14716 32635
rect 14531 32585 14606 32601
rect 14640 32585 14716 32619
rect 14531 32567 14716 32585
rect 14531 32533 14599 32567
rect 14633 32547 14716 32567
rect 14531 32513 14606 32533
rect 14640 32513 14716 32547
rect 14531 32499 14716 32513
rect 14531 32465 14599 32499
rect 14633 32475 14716 32499
rect 14531 32441 14606 32465
rect 14640 32441 14716 32475
rect 14531 32431 14716 32441
rect 14531 32397 14599 32431
rect 14633 32403 14716 32431
rect 14531 32369 14606 32397
rect 14640 32369 14716 32403
rect 14531 32363 14716 32369
rect 14531 32329 14599 32363
rect 14633 32331 14716 32363
rect 14531 32297 14606 32329
rect 14640 32297 14716 32331
rect 14531 32295 14716 32297
rect 14531 32261 14599 32295
rect 14633 32261 14716 32295
rect 14531 32259 14716 32261
rect 14531 32227 14606 32259
rect 14531 32193 14599 32227
rect 14640 32225 14716 32259
rect 14633 32193 14716 32225
rect 14531 32187 14716 32193
rect 14531 32159 14606 32187
rect 14531 32125 14599 32159
rect 14640 32153 14716 32187
rect 14633 32125 14716 32153
rect 14531 32115 14716 32125
rect 14531 32091 14606 32115
rect 14531 32057 14599 32091
rect 14640 32081 14716 32115
rect 14633 32057 14716 32081
rect 14531 32043 14716 32057
rect 14531 32023 14606 32043
rect 14531 31989 14599 32023
rect 14640 32009 14716 32043
rect 14633 31989 14716 32009
rect 14531 31971 14716 31989
rect 14531 31955 14606 31971
rect 14531 31921 14599 31955
rect 14640 31937 14716 31971
rect 14633 31921 14716 31937
rect 14531 31899 14716 31921
rect 14531 31887 14606 31899
rect 14531 31853 14599 31887
rect 14640 31865 14716 31899
rect 14633 31853 14716 31865
rect 14531 31827 14716 31853
rect 14531 31819 14606 31827
rect 14531 31785 14599 31819
rect 14640 31793 14716 31827
rect 14633 31785 14716 31793
rect 14531 31755 14716 31785
rect 14531 31751 14606 31755
rect 14531 31717 14599 31751
rect 14640 31721 14716 31755
rect 14633 31717 14716 31721
rect 14531 31683 14716 31717
rect 14531 31649 14599 31683
rect 14640 31649 14716 31683
rect 14531 31615 14716 31649
rect 14531 31581 14599 31615
rect 14633 31611 14716 31615
rect 14531 31577 14606 31581
rect 14640 31577 14716 31611
rect 14531 31547 14716 31577
rect 14531 31513 14599 31547
rect 14633 31539 14716 31547
rect 14531 31505 14606 31513
rect 14640 31505 14716 31539
rect 14531 31479 14716 31505
rect 14531 31445 14599 31479
rect 14633 31467 14716 31479
rect 14531 31433 14606 31445
rect 14640 31433 14716 31467
rect 14531 31411 14716 31433
rect 14531 31377 14599 31411
rect 14633 31395 14716 31411
rect 14531 31361 14606 31377
rect 14640 31361 14716 31395
rect 14531 31343 14716 31361
rect 14531 31309 14599 31343
rect 14633 31323 14716 31343
rect 14531 31289 14606 31309
rect 14640 31289 14716 31323
rect 14531 31275 14716 31289
rect 14531 31241 14599 31275
rect 14633 31251 14716 31275
rect 14531 31217 14606 31241
rect 14640 31217 14716 31251
rect 14531 31207 14716 31217
rect 14531 31173 14599 31207
rect 14633 31179 14716 31207
rect 14531 31145 14606 31173
rect 14640 31145 14716 31179
rect 14531 31139 14716 31145
rect 14531 31105 14599 31139
rect 14633 31107 14716 31139
rect 14531 31073 14606 31105
rect 14640 31073 14716 31107
rect 14531 31071 14716 31073
rect 14531 31037 14599 31071
rect 14633 31037 14716 31071
rect 14531 31035 14716 31037
rect 14531 31003 14606 31035
rect 14531 30969 14599 31003
rect 14640 31001 14716 31035
rect 14633 30969 14716 31001
rect 14531 30963 14716 30969
rect 14531 30935 14606 30963
rect 14531 30901 14599 30935
rect 14640 30929 14716 30963
rect 14633 30901 14716 30929
rect 14531 30891 14716 30901
rect 14531 30867 14606 30891
rect 14531 30833 14599 30867
rect 14640 30857 14716 30891
rect 14633 30833 14716 30857
rect 14531 30819 14716 30833
rect 14531 30799 14606 30819
rect 14531 30765 14599 30799
rect 14640 30785 14716 30819
rect 14633 30765 14716 30785
rect 14531 30747 14716 30765
rect 14531 30731 14606 30747
rect 14531 30697 14599 30731
rect 14640 30713 14716 30747
rect 14633 30697 14716 30713
rect 14531 30675 14716 30697
rect 14531 30663 14606 30675
rect 14531 30629 14599 30663
rect 14640 30641 14716 30675
rect 14633 30629 14716 30641
rect 14531 30603 14716 30629
rect 14531 30595 14606 30603
rect 14531 30561 14599 30595
rect 14640 30569 14716 30603
rect 14633 30561 14716 30569
rect 14531 30531 14716 30561
rect 14531 30527 14606 30531
rect 14531 30493 14599 30527
rect 14640 30497 14716 30531
rect 14633 30493 14716 30497
rect 14531 30459 14716 30493
rect 14531 30425 14599 30459
rect 14640 30425 14716 30459
rect 14531 30391 14716 30425
rect 14531 30357 14599 30391
rect 14633 30387 14716 30391
rect 14531 30353 14606 30357
rect 14640 30353 14716 30387
rect 14531 30323 14716 30353
rect 14531 30289 14599 30323
rect 14633 30315 14716 30323
rect 14531 30281 14606 30289
rect 14640 30281 14716 30315
rect 14531 30255 14716 30281
rect 14531 30221 14599 30255
rect 14633 30243 14716 30255
rect 14531 30209 14606 30221
rect 14640 30209 14716 30243
rect 14531 30187 14716 30209
rect 14531 30153 14599 30187
rect 14633 30171 14716 30187
rect 14531 30137 14606 30153
rect 14640 30137 14716 30171
rect 14531 30119 14716 30137
rect 14531 30085 14599 30119
rect 14633 30099 14716 30119
rect 14531 30065 14606 30085
rect 14640 30065 14716 30099
rect 14531 30051 14716 30065
rect 14531 30017 14599 30051
rect 14633 30027 14716 30051
rect 14531 29993 14606 30017
rect 14640 29993 14716 30027
rect 14531 29983 14716 29993
rect 14531 29949 14599 29983
rect 14633 29955 14716 29983
rect 14531 29921 14606 29949
rect 14640 29921 14716 29955
rect 14531 29915 14716 29921
rect 14531 29881 14599 29915
rect 14633 29883 14716 29915
rect 14531 29849 14606 29881
rect 14640 29849 14716 29883
rect 14531 29847 14716 29849
rect 14531 29813 14599 29847
rect 14633 29813 14716 29847
rect 14531 29811 14716 29813
rect 14531 29779 14606 29811
rect 14531 29745 14599 29779
rect 14640 29777 14716 29811
rect 14633 29745 14716 29777
rect 14531 29739 14716 29745
rect 14531 29711 14606 29739
rect 14531 29677 14599 29711
rect 14640 29705 14716 29739
rect 14633 29677 14716 29705
rect 14531 29667 14716 29677
rect 14531 29643 14606 29667
rect 14531 29609 14599 29643
rect 14640 29633 14716 29667
rect 14633 29609 14716 29633
rect 14531 29595 14716 29609
rect 14531 29575 14606 29595
rect 14531 29541 14599 29575
rect 14640 29561 14716 29595
rect 14633 29541 14716 29561
rect 14531 29523 14716 29541
rect 14531 29507 14606 29523
rect 14531 29473 14599 29507
rect 14640 29489 14716 29523
rect 14633 29473 14716 29489
rect 14531 29451 14716 29473
rect 14531 29439 14606 29451
rect 14531 29405 14599 29439
rect 14640 29417 14716 29451
rect 14633 29405 14716 29417
rect 14531 29379 14716 29405
rect 14531 29371 14606 29379
rect 14531 29337 14599 29371
rect 14640 29345 14716 29379
rect 14633 29337 14716 29345
rect 14531 29307 14716 29337
rect 14531 29303 14606 29307
rect 14531 29269 14599 29303
rect 14640 29273 14716 29307
rect 14633 29269 14716 29273
rect 14531 29235 14716 29269
rect 14531 29201 14599 29235
rect 14640 29201 14716 29235
rect 14531 29167 14716 29201
rect 14531 29133 14599 29167
rect 14633 29163 14716 29167
rect 14531 29129 14606 29133
rect 14640 29129 14716 29163
rect 14531 29099 14716 29129
rect 14531 29065 14599 29099
rect 14633 29091 14716 29099
rect 14531 29057 14606 29065
rect 14640 29057 14716 29091
rect 14531 29031 14716 29057
rect 14531 28997 14599 29031
rect 14633 29019 14716 29031
rect 14531 28985 14606 28997
rect 14640 28985 14716 29019
rect 14531 28963 14716 28985
rect 14531 28929 14599 28963
rect 14633 28947 14716 28963
rect 14531 28913 14606 28929
rect 14640 28913 14716 28947
rect 14531 28895 14716 28913
rect 14531 28861 14599 28895
rect 14633 28875 14716 28895
rect 14531 28841 14606 28861
rect 14640 28841 14716 28875
rect 14531 28827 14716 28841
rect 14531 28793 14599 28827
rect 14633 28803 14716 28827
rect 14531 28769 14606 28793
rect 14640 28769 14716 28803
rect 14531 28759 14716 28769
rect 14531 28725 14599 28759
rect 14633 28731 14716 28759
rect 14531 28697 14606 28725
rect 14640 28697 14716 28731
rect 14531 28691 14716 28697
rect 14531 28657 14599 28691
rect 14633 28659 14716 28691
rect 14531 28625 14606 28657
rect 14640 28625 14716 28659
rect 14531 28623 14716 28625
rect 14531 28589 14599 28623
rect 14633 28589 14716 28623
rect 14531 28587 14716 28589
rect 14531 28555 14606 28587
rect 14531 28521 14599 28555
rect 14640 28553 14716 28587
rect 14633 28521 14716 28553
rect 14531 28515 14716 28521
rect 14531 28487 14606 28515
rect 14531 28453 14599 28487
rect 14640 28481 14716 28515
rect 14633 28453 14716 28481
rect 14531 28443 14716 28453
rect 14531 28419 14606 28443
rect 14531 28385 14599 28419
rect 14640 28409 14716 28443
rect 14633 28385 14716 28409
rect 14531 28371 14716 28385
rect 14531 28351 14606 28371
rect 14531 28317 14599 28351
rect 14640 28337 14716 28371
rect 14633 28317 14716 28337
rect 14531 28299 14716 28317
rect 14531 28283 14606 28299
rect 14531 28249 14599 28283
rect 14640 28265 14716 28299
rect 14633 28249 14716 28265
rect 14531 28227 14716 28249
rect 14531 28215 14606 28227
rect 14531 28181 14599 28215
rect 14640 28193 14716 28227
rect 14633 28181 14716 28193
rect 14531 28155 14716 28181
rect 14531 28147 14606 28155
rect 14531 28113 14599 28147
rect 14640 28121 14716 28155
rect 14633 28113 14716 28121
rect 14531 28083 14716 28113
rect 14531 28079 14606 28083
rect 14531 28045 14599 28079
rect 14640 28049 14716 28083
rect 14633 28045 14716 28049
rect 14531 28011 14716 28045
rect 14531 27977 14599 28011
rect 14640 27977 14716 28011
rect 14531 27943 14716 27977
rect 14531 27909 14599 27943
rect 14633 27939 14716 27943
rect 14531 27905 14606 27909
rect 14640 27905 14716 27939
rect 14531 27875 14716 27905
rect 14531 27841 14599 27875
rect 14633 27867 14716 27875
rect 14531 27833 14606 27841
rect 14640 27833 14716 27867
rect 14531 27807 14716 27833
rect 14531 27773 14599 27807
rect 14633 27795 14716 27807
rect 14531 27761 14606 27773
rect 14640 27761 14716 27795
rect 14531 27739 14716 27761
rect 14531 27705 14599 27739
rect 14633 27723 14716 27739
rect 14531 27689 14606 27705
rect 14640 27689 14716 27723
rect 14531 27671 14716 27689
rect 14531 27637 14599 27671
rect 14633 27651 14716 27671
rect 14531 27617 14606 27637
rect 14640 27617 14716 27651
rect 14531 27603 14716 27617
rect 14531 27569 14599 27603
rect 14633 27579 14716 27603
rect 14531 27545 14606 27569
rect 14640 27545 14716 27579
rect 14531 27535 14716 27545
rect 14531 27501 14599 27535
rect 14633 27507 14716 27535
rect 14531 27473 14606 27501
rect 14640 27473 14716 27507
rect 14531 27467 14716 27473
rect 14531 27433 14599 27467
rect 14633 27435 14716 27467
rect 14531 27401 14606 27433
rect 14640 27401 14716 27435
rect 14531 27399 14716 27401
rect 14531 27365 14599 27399
rect 14633 27365 14716 27399
rect 14531 27363 14716 27365
rect 14531 27331 14606 27363
rect 14531 27297 14599 27331
rect 14640 27329 14716 27363
rect 14633 27297 14716 27329
rect 14531 27291 14716 27297
rect 14531 27263 14606 27291
rect 14531 27229 14599 27263
rect 14640 27257 14716 27291
rect 14633 27229 14716 27257
rect 14531 27219 14716 27229
rect 14531 27195 14606 27219
rect 14531 27161 14599 27195
rect 14640 27185 14716 27219
rect 14633 27161 14716 27185
rect 14531 27147 14716 27161
rect 14531 27127 14606 27147
rect 14531 27093 14599 27127
rect 14640 27113 14716 27147
rect 14633 27093 14716 27113
rect 14531 27075 14716 27093
rect 14531 27059 14606 27075
rect 14531 27025 14599 27059
rect 14640 27041 14716 27075
rect 14633 27025 14716 27041
rect 14531 27003 14716 27025
rect 14531 26991 14606 27003
rect 14531 26957 14599 26991
rect 14640 26969 14716 27003
rect 14633 26957 14716 26969
rect 14531 26931 14716 26957
rect 14531 26923 14606 26931
rect 14531 26889 14599 26923
rect 14640 26897 14716 26931
rect 14633 26889 14716 26897
rect 14531 26859 14716 26889
rect 14531 26855 14606 26859
rect 14531 26821 14599 26855
rect 14640 26825 14716 26859
rect 14633 26821 14716 26825
rect 14531 26787 14716 26821
rect 14531 26753 14599 26787
rect 14640 26753 14716 26787
rect 14531 26719 14716 26753
rect 14531 26685 14599 26719
rect 14633 26715 14716 26719
rect 14531 26681 14606 26685
rect 14640 26681 14716 26715
rect 14531 26651 14716 26681
rect 14531 26617 14599 26651
rect 14633 26643 14716 26651
rect 14531 26609 14606 26617
rect 14640 26609 14716 26643
rect 14531 26583 14716 26609
rect 14531 26549 14599 26583
rect 14633 26571 14716 26583
rect 14531 26537 14606 26549
rect 14640 26537 14716 26571
rect 14531 26515 14716 26537
rect 14531 26481 14599 26515
rect 14633 26499 14716 26515
rect 14531 26465 14606 26481
rect 14640 26465 14716 26499
rect 14531 26447 14716 26465
rect 14531 26413 14599 26447
rect 14633 26427 14716 26447
rect 14531 26393 14606 26413
rect 14640 26393 14716 26427
rect 14531 26379 14716 26393
rect 14531 26345 14599 26379
rect 14633 26355 14716 26379
rect 14531 26321 14606 26345
rect 14640 26321 14716 26355
rect 14531 26311 14716 26321
rect 14531 26277 14599 26311
rect 14633 26283 14716 26311
rect 14531 26249 14606 26277
rect 14640 26249 14716 26283
rect 14531 26243 14716 26249
rect 14531 26209 14599 26243
rect 14633 26211 14716 26243
rect 14531 26177 14606 26209
rect 14640 26177 14716 26211
rect 14531 26175 14716 26177
rect 14531 26141 14599 26175
rect 14633 26141 14716 26175
rect 14531 26139 14716 26141
rect 14531 26107 14606 26139
rect 14531 26073 14599 26107
rect 14640 26105 14716 26139
rect 14633 26073 14716 26105
rect 14531 26067 14716 26073
rect 14531 26039 14606 26067
rect 14531 26005 14599 26039
rect 14640 26033 14716 26067
rect 14633 26005 14716 26033
rect 14531 25995 14716 26005
rect 14531 25971 14606 25995
rect 14531 25937 14599 25971
rect 14640 25961 14716 25995
rect 14633 25937 14716 25961
rect 14531 25923 14716 25937
rect 14531 25903 14606 25923
rect 14531 25869 14599 25903
rect 14640 25889 14716 25923
rect 14633 25869 14716 25889
rect 14531 25851 14716 25869
rect 14531 25835 14606 25851
rect 14531 25801 14599 25835
rect 14640 25817 14716 25851
rect 14633 25801 14716 25817
rect 14531 25779 14716 25801
rect 14531 25767 14606 25779
rect 14531 25733 14599 25767
rect 14640 25745 14716 25779
rect 14633 25733 14716 25745
rect 14531 25707 14716 25733
rect 14531 25699 14606 25707
rect 14531 25665 14599 25699
rect 14640 25673 14716 25707
rect 14633 25665 14716 25673
rect 14531 25635 14716 25665
rect 14531 25631 14606 25635
rect 14531 25597 14599 25631
rect 14640 25601 14716 25635
rect 14633 25597 14716 25601
rect 14531 25563 14716 25597
rect 14531 25529 14599 25563
rect 14640 25529 14716 25563
rect 14531 25495 14716 25529
rect 14531 25461 14599 25495
rect 14633 25491 14716 25495
rect 14531 25457 14606 25461
rect 14640 25457 14716 25491
rect 14531 25427 14716 25457
rect 14531 25393 14599 25427
rect 14633 25419 14716 25427
rect 14531 25385 14606 25393
rect 14640 25385 14716 25419
rect 14531 25359 14716 25385
rect 14531 25325 14599 25359
rect 14633 25347 14716 25359
rect 14531 25313 14606 25325
rect 14640 25313 14716 25347
rect 14531 25291 14716 25313
rect 14531 25257 14599 25291
rect 14633 25275 14716 25291
rect 14531 25241 14606 25257
rect 14640 25241 14716 25275
rect 14531 25223 14716 25241
rect 14531 25189 14599 25223
rect 14633 25203 14716 25223
rect 14531 25169 14606 25189
rect 14640 25169 14716 25203
rect 14531 25155 14716 25169
rect 14531 25121 14599 25155
rect 14633 25131 14716 25155
rect 14531 25097 14606 25121
rect 14640 25097 14716 25131
rect 14531 25087 14716 25097
rect 14531 25053 14599 25087
rect 14633 25059 14716 25087
rect 14531 25025 14606 25053
rect 14640 25025 14716 25059
rect 14531 25019 14716 25025
rect 14531 24985 14599 25019
rect 14633 24987 14716 25019
rect 14531 24953 14606 24985
rect 14640 24953 14716 24987
rect 14531 24951 14716 24953
rect 14531 24917 14599 24951
rect 14633 24917 14716 24951
rect 14531 24915 14716 24917
rect 14531 24883 14606 24915
rect 14531 24849 14599 24883
rect 14640 24881 14716 24915
rect 14633 24849 14716 24881
rect 14531 24843 14716 24849
rect 14531 24815 14606 24843
rect 14531 24781 14599 24815
rect 14640 24809 14716 24843
rect 14633 24781 14716 24809
rect 14531 24771 14716 24781
rect 14531 24747 14606 24771
rect 14531 24713 14599 24747
rect 14640 24737 14716 24771
rect 14633 24713 14716 24737
rect 14531 24699 14716 24713
rect 14531 24679 14606 24699
rect 14531 24645 14599 24679
rect 14640 24665 14716 24699
rect 14633 24645 14716 24665
rect 14531 24627 14716 24645
rect 14531 24611 14606 24627
rect 14531 24577 14599 24611
rect 14640 24593 14716 24627
rect 14633 24577 14716 24593
rect 14531 24555 14716 24577
rect 14531 24543 14606 24555
rect 14531 24509 14599 24543
rect 14640 24521 14716 24555
rect 14633 24509 14716 24521
rect 14531 24483 14716 24509
rect 14531 24475 14606 24483
rect 14531 24441 14599 24475
rect 14640 24449 14716 24483
rect 14633 24441 14716 24449
rect 14531 24411 14716 24441
rect 14531 24407 14606 24411
rect 14531 24373 14599 24407
rect 14640 24377 14716 24411
rect 14633 24373 14716 24377
rect 14531 24339 14716 24373
rect 14531 24305 14599 24339
rect 14640 24305 14716 24339
rect 14531 24271 14716 24305
rect 14531 24237 14599 24271
rect 14633 24267 14716 24271
rect 14531 24233 14606 24237
rect 14640 24233 14716 24267
rect 14531 24203 14716 24233
rect 14531 24169 14599 24203
rect 14633 24195 14716 24203
rect 14531 24161 14606 24169
rect 14640 24161 14716 24195
rect 14531 24135 14716 24161
rect 14531 24101 14599 24135
rect 14633 24123 14716 24135
rect 14531 24089 14606 24101
rect 14640 24089 14716 24123
rect 14531 24067 14716 24089
rect 14531 24033 14599 24067
rect 14633 24051 14716 24067
rect 14531 24017 14606 24033
rect 14640 24017 14716 24051
rect 14531 23999 14716 24017
rect 14531 23965 14599 23999
rect 14633 23979 14716 23999
rect 14531 23945 14606 23965
rect 14640 23945 14716 23979
rect 14531 23931 14716 23945
rect 14531 23897 14599 23931
rect 14633 23907 14716 23931
rect 14531 23873 14606 23897
rect 14640 23873 14716 23907
rect 14531 23863 14716 23873
rect 14531 23829 14599 23863
rect 14633 23835 14716 23863
rect 14531 23801 14606 23829
rect 14640 23801 14716 23835
rect 14531 23795 14716 23801
rect 14531 23761 14599 23795
rect 14633 23763 14716 23795
rect 14531 23729 14606 23761
rect 14640 23729 14716 23763
rect 14531 23727 14716 23729
rect 14531 23693 14599 23727
rect 14633 23693 14716 23727
rect 14531 23691 14716 23693
rect 14531 23659 14606 23691
rect 14531 23625 14599 23659
rect 14640 23657 14716 23691
rect 14633 23625 14716 23657
rect 14531 23619 14716 23625
rect 14531 23591 14606 23619
rect 14531 23557 14599 23591
rect 14640 23585 14716 23619
rect 14633 23557 14716 23585
rect 14531 23547 14716 23557
rect 14531 23523 14606 23547
rect 14531 23489 14599 23523
rect 14640 23513 14716 23547
rect 14633 23489 14716 23513
rect 14531 23475 14716 23489
rect 14531 23455 14606 23475
rect 14531 23421 14599 23455
rect 14640 23441 14716 23475
rect 14633 23421 14716 23441
rect 14531 23403 14716 23421
rect 14531 23387 14606 23403
rect 14531 23353 14599 23387
rect 14640 23369 14716 23403
rect 14633 23353 14716 23369
rect 14531 23331 14716 23353
rect 14531 23319 14606 23331
rect 14531 23285 14599 23319
rect 14640 23297 14716 23331
rect 14633 23285 14716 23297
rect 14531 23259 14716 23285
rect 14531 23251 14606 23259
rect 14531 23217 14599 23251
rect 14640 23225 14716 23259
rect 14633 23217 14716 23225
rect 14531 23187 14716 23217
rect 14531 23183 14606 23187
rect 14531 23149 14599 23183
rect 14640 23153 14716 23187
rect 14633 23149 14716 23153
rect 14531 23115 14716 23149
rect 14531 23081 14599 23115
rect 14640 23081 14716 23115
rect 14531 23047 14716 23081
rect 14531 23013 14599 23047
rect 14633 23043 14716 23047
rect 14531 23009 14606 23013
rect 14640 23009 14716 23043
rect 14531 22979 14716 23009
rect 14531 22945 14599 22979
rect 14633 22971 14716 22979
rect 14531 22937 14606 22945
rect 14640 22937 14716 22971
rect 14531 22911 14716 22937
rect 14531 22877 14599 22911
rect 14633 22899 14716 22911
rect 14531 22865 14606 22877
rect 14640 22865 14716 22899
rect 14531 22843 14716 22865
rect 14531 22809 14599 22843
rect 14633 22827 14716 22843
rect 14531 22793 14606 22809
rect 14640 22793 14716 22827
rect 14531 22775 14716 22793
rect 14531 22741 14599 22775
rect 14633 22755 14716 22775
rect 14531 22721 14606 22741
rect 14640 22721 14716 22755
rect 14531 22707 14716 22721
rect 14531 22673 14599 22707
rect 14633 22683 14716 22707
rect 14531 22649 14606 22673
rect 14640 22649 14716 22683
rect 14531 22639 14716 22649
rect 14531 22605 14599 22639
rect 14633 22611 14716 22639
rect 14531 22577 14606 22605
rect 14640 22577 14716 22611
rect 14531 22571 14716 22577
rect 14531 22537 14599 22571
rect 14633 22539 14716 22571
rect 14531 22505 14606 22537
rect 14640 22505 14716 22539
rect 14531 22503 14716 22505
rect 14531 22469 14599 22503
rect 14633 22469 14716 22503
rect 14531 22467 14716 22469
rect 14531 22435 14606 22467
rect 14531 22401 14599 22435
rect 14640 22433 14716 22467
rect 14633 22401 14716 22433
rect 14531 22395 14716 22401
rect 14531 22367 14606 22395
rect 14531 22333 14599 22367
rect 14640 22361 14716 22395
rect 14633 22333 14716 22361
rect 14531 22323 14716 22333
rect 14531 22299 14606 22323
rect 14531 22265 14599 22299
rect 14640 22289 14716 22323
rect 14633 22265 14716 22289
rect 14531 22251 14716 22265
rect 14531 22231 14606 22251
rect 14531 22197 14599 22231
rect 14640 22217 14716 22251
rect 14633 22197 14716 22217
rect 14531 22179 14716 22197
rect 14531 22163 14606 22179
rect 14531 22129 14599 22163
rect 14640 22145 14716 22179
rect 14633 22129 14716 22145
rect 14531 22107 14716 22129
rect 14531 22095 14606 22107
rect 14531 22061 14599 22095
rect 14640 22073 14716 22107
rect 14633 22061 14716 22073
rect 14531 22035 14716 22061
rect 14531 22027 14606 22035
rect 14531 21993 14599 22027
rect 14640 22001 14716 22035
rect 14633 21993 14716 22001
rect 14531 21963 14716 21993
rect 14531 21959 14606 21963
rect 14531 21925 14599 21959
rect 14640 21929 14716 21963
rect 14633 21925 14716 21929
rect 14531 21891 14716 21925
rect 14531 21857 14599 21891
rect 14640 21857 14716 21891
rect 14531 21823 14716 21857
rect 14531 21789 14599 21823
rect 14633 21819 14716 21823
rect 14531 21785 14606 21789
rect 14640 21785 14716 21819
rect 14531 21755 14716 21785
rect 14531 21721 14599 21755
rect 14633 21747 14716 21755
rect 14531 21713 14606 21721
rect 14640 21713 14716 21747
rect 14531 21687 14716 21713
rect 14531 21653 14599 21687
rect 14633 21675 14716 21687
rect 14531 21641 14606 21653
rect 14640 21641 14716 21675
rect 14531 21619 14716 21641
rect 14531 21585 14599 21619
rect 14633 21603 14716 21619
rect 14531 21569 14606 21585
rect 14640 21569 14716 21603
rect 14531 21551 14716 21569
rect 14531 21517 14599 21551
rect 14633 21531 14716 21551
rect 14531 21497 14606 21517
rect 14640 21497 14716 21531
rect 14531 21483 14716 21497
rect 14531 21449 14599 21483
rect 14633 21459 14716 21483
rect 14531 21425 14606 21449
rect 14640 21425 14716 21459
rect 14531 21415 14716 21425
rect 14531 21381 14599 21415
rect 14633 21387 14716 21415
rect 14531 21353 14606 21381
rect 14640 21353 14716 21387
rect 14531 21347 14716 21353
rect 14531 21313 14599 21347
rect 14633 21315 14716 21347
rect 14531 21281 14606 21313
rect 14640 21281 14716 21315
rect 14531 21279 14716 21281
rect 14531 21245 14599 21279
rect 14633 21245 14716 21279
rect 14531 21243 14716 21245
rect 14531 21211 14606 21243
rect 14531 21177 14599 21211
rect 14640 21209 14716 21243
rect 14633 21177 14716 21209
rect 14531 21171 14716 21177
rect 14531 21143 14606 21171
rect 14531 21109 14599 21143
rect 14640 21137 14716 21171
rect 14633 21109 14716 21137
rect 14531 21099 14716 21109
rect 14531 21075 14606 21099
rect 14531 21041 14599 21075
rect 14640 21065 14716 21099
rect 14633 21041 14716 21065
rect 14531 21027 14716 21041
rect 14531 21007 14606 21027
rect 14531 20973 14599 21007
rect 14640 20993 14716 21027
rect 14633 20973 14716 20993
rect 14531 20955 14716 20973
rect 14531 20939 14606 20955
rect 14531 20905 14599 20939
rect 14640 20921 14716 20955
rect 14633 20905 14716 20921
rect 14531 20883 14716 20905
rect 14531 20871 14606 20883
rect 14531 20837 14599 20871
rect 14640 20849 14716 20883
rect 14633 20837 14716 20849
rect 14531 20811 14716 20837
rect 14531 20803 14606 20811
rect 14531 20769 14599 20803
rect 14640 20777 14716 20811
rect 14633 20769 14716 20777
rect 14531 20739 14716 20769
rect 14531 20735 14606 20739
rect 14531 20701 14599 20735
rect 14640 20705 14716 20739
rect 14633 20701 14716 20705
rect 14531 20667 14716 20701
rect 14531 20633 14599 20667
rect 14640 20633 14716 20667
rect 14531 20599 14716 20633
rect 14531 20565 14599 20599
rect 14633 20595 14716 20599
rect 14531 20561 14606 20565
rect 14640 20561 14716 20595
rect 14531 20531 14716 20561
rect 14531 20497 14599 20531
rect 14633 20523 14716 20531
rect 14531 20489 14606 20497
rect 14640 20489 14716 20523
rect 14531 20463 14716 20489
rect 14531 20429 14599 20463
rect 14633 20451 14716 20463
rect 14531 20417 14606 20429
rect 14640 20417 14716 20451
rect 14531 20395 14716 20417
rect 14531 20361 14599 20395
rect 14633 20379 14716 20395
rect 14531 20345 14606 20361
rect 14640 20345 14716 20379
rect 14531 20327 14716 20345
rect 14531 20293 14599 20327
rect 14633 20307 14716 20327
rect 14531 20273 14606 20293
rect 14640 20273 14716 20307
rect 14531 20259 14716 20273
rect 14531 20225 14599 20259
rect 14633 20235 14716 20259
rect 14531 20201 14606 20225
rect 14640 20201 14716 20235
rect 14531 20191 14716 20201
rect 14531 20157 14599 20191
rect 14633 20163 14716 20191
rect 14531 20129 14606 20157
rect 14640 20129 14716 20163
rect 14531 20123 14716 20129
rect 14531 20089 14599 20123
rect 14633 20091 14716 20123
rect 14531 20057 14606 20089
rect 14640 20057 14716 20091
rect 14531 20055 14716 20057
rect 14531 20021 14599 20055
rect 14633 20021 14716 20055
rect 14531 20019 14716 20021
rect 14531 19987 14606 20019
rect 14531 19953 14599 19987
rect 14640 19985 14716 20019
rect 14633 19953 14716 19985
rect 14531 19947 14716 19953
rect 14531 19919 14606 19947
rect 14531 19885 14599 19919
rect 14640 19913 14716 19947
rect 14633 19885 14716 19913
rect 14531 19875 14716 19885
rect 14531 19851 14606 19875
rect 14531 19817 14599 19851
rect 14640 19841 14716 19875
rect 14633 19817 14716 19841
rect 14531 19803 14716 19817
rect 14531 19783 14606 19803
rect 14531 19749 14599 19783
rect 14640 19769 14716 19803
rect 14633 19749 14716 19769
rect 14531 19731 14716 19749
rect 14531 19715 14606 19731
rect 14531 19681 14599 19715
rect 14640 19697 14716 19731
rect 14633 19681 14716 19697
rect 14531 19659 14716 19681
rect 14531 19647 14606 19659
rect 14531 19613 14599 19647
rect 14640 19625 14716 19659
rect 14633 19613 14716 19625
rect 14531 19587 14716 19613
rect 14531 19579 14606 19587
rect 14531 19545 14599 19579
rect 14640 19553 14716 19587
rect 14633 19545 14716 19553
rect 14531 19515 14716 19545
rect 14531 19511 14606 19515
rect 14531 19477 14599 19511
rect 14640 19481 14716 19515
rect 14633 19477 14716 19481
rect 14531 19443 14716 19477
rect 14531 19409 14599 19443
rect 14640 19409 14716 19443
rect 14531 19375 14716 19409
rect 14531 19341 14599 19375
rect 14633 19371 14716 19375
rect 14531 19337 14606 19341
rect 14640 19337 14716 19371
rect 14531 19307 14716 19337
rect 14531 19273 14599 19307
rect 14633 19299 14716 19307
rect 14531 19265 14606 19273
rect 14640 19265 14716 19299
rect 14531 19239 14716 19265
rect 14531 19205 14599 19239
rect 14633 19227 14716 19239
rect 14531 19193 14606 19205
rect 14640 19193 14716 19227
rect 14531 19171 14716 19193
rect 14531 19137 14599 19171
rect 14633 19155 14716 19171
rect 14531 19121 14606 19137
rect 14640 19121 14716 19155
rect 14531 19103 14716 19121
rect 14531 19069 14599 19103
rect 14633 19083 14716 19103
rect 14531 19049 14606 19069
rect 14640 19049 14716 19083
rect 14531 19035 14716 19049
rect 14531 19001 14599 19035
rect 14633 19011 14716 19035
rect 14531 18977 14606 19001
rect 14640 18977 14716 19011
rect 14531 18967 14716 18977
rect 14531 18933 14599 18967
rect 14633 18939 14716 18967
rect 14531 18905 14606 18933
rect 14640 18905 14716 18939
rect 14531 18899 14716 18905
rect 14531 18865 14599 18899
rect 14633 18867 14716 18899
rect 14531 18833 14606 18865
rect 14640 18833 14716 18867
rect 14531 18831 14716 18833
rect 14531 18797 14599 18831
rect 14633 18797 14716 18831
rect 14531 18795 14716 18797
rect 14531 18763 14606 18795
rect 14531 18729 14599 18763
rect 14640 18761 14716 18795
rect 14633 18729 14716 18761
rect 14531 18723 14716 18729
rect 14531 18695 14606 18723
rect 14531 18661 14599 18695
rect 14640 18689 14716 18723
rect 14633 18661 14716 18689
rect 14531 18651 14716 18661
rect 14531 18627 14606 18651
rect 14531 18593 14599 18627
rect 14640 18617 14716 18651
rect 14633 18593 14716 18617
rect 14531 18579 14716 18593
rect 14531 18559 14606 18579
rect 14531 18525 14599 18559
rect 14640 18545 14716 18579
rect 14633 18525 14716 18545
rect 14531 18507 14716 18525
rect 14531 18491 14606 18507
rect 14531 18457 14599 18491
rect 14640 18473 14716 18507
rect 14633 18457 14716 18473
rect 14531 18435 14716 18457
rect 14531 18423 14606 18435
rect 14531 18389 14599 18423
rect 14640 18401 14716 18435
rect 14633 18389 14716 18401
rect 14531 18363 14716 18389
rect 14531 18355 14606 18363
rect 14531 18321 14599 18355
rect 14640 18329 14716 18363
rect 14633 18321 14716 18329
rect 14531 18291 14716 18321
rect 14531 18287 14606 18291
rect 14531 18253 14599 18287
rect 14640 18257 14716 18291
rect 14633 18253 14716 18257
rect 14531 18219 14716 18253
rect 14531 18185 14599 18219
rect 14640 18185 14716 18219
rect 14531 18151 14716 18185
rect 14531 18117 14599 18151
rect 14633 18147 14716 18151
rect 14531 18113 14606 18117
rect 14640 18113 14716 18147
rect 14531 18083 14716 18113
rect 14531 18049 14599 18083
rect 14633 18075 14716 18083
rect 14531 18041 14606 18049
rect 14640 18041 14716 18075
rect 14531 18015 14716 18041
rect 14531 17981 14599 18015
rect 14633 18003 14716 18015
rect 14531 17969 14606 17981
rect 14640 17969 14716 18003
rect 14531 17947 14716 17969
rect 14531 17913 14599 17947
rect 14633 17931 14716 17947
rect 14531 17897 14606 17913
rect 14640 17897 14716 17931
rect 14531 17879 14716 17897
rect 14531 17845 14599 17879
rect 14633 17859 14716 17879
rect 14531 17825 14606 17845
rect 14640 17825 14716 17859
rect 14531 17811 14716 17825
rect 14531 17777 14599 17811
rect 14633 17787 14716 17811
rect 14531 17753 14606 17777
rect 14640 17753 14716 17787
rect 14531 17743 14716 17753
rect 14531 17709 14599 17743
rect 14633 17715 14716 17743
rect 14531 17681 14606 17709
rect 14640 17681 14716 17715
rect 14531 17675 14716 17681
rect 14531 17641 14599 17675
rect 14633 17643 14716 17675
rect 14531 17609 14606 17641
rect 14640 17609 14716 17643
rect 14531 17607 14716 17609
rect 14531 17573 14599 17607
rect 14633 17573 14716 17607
rect 14531 17571 14716 17573
rect 14531 17539 14606 17571
rect 14531 17505 14599 17539
rect 14640 17537 14716 17571
rect 14633 17505 14716 17537
rect 14531 17499 14716 17505
rect 14531 17471 14606 17499
rect 14531 17437 14599 17471
rect 14640 17465 14716 17499
rect 14633 17437 14716 17465
rect 14531 17427 14716 17437
rect 14531 17403 14606 17427
rect 14531 17369 14599 17403
rect 14640 17393 14716 17427
rect 14633 17369 14716 17393
rect 14531 17355 14716 17369
rect 14531 17335 14606 17355
rect 14531 17301 14599 17335
rect 14640 17321 14716 17355
rect 14633 17301 14716 17321
rect 14531 17283 14716 17301
rect 14531 17267 14606 17283
rect 14531 17233 14599 17267
rect 14640 17249 14716 17283
rect 14633 17233 14716 17249
rect 14531 17211 14716 17233
rect 14531 17199 14606 17211
rect 14531 17165 14599 17199
rect 14640 17177 14716 17211
rect 14633 17165 14716 17177
rect 14531 17139 14716 17165
rect 14531 17131 14606 17139
rect 14531 17097 14599 17131
rect 14640 17105 14716 17139
rect 14633 17097 14716 17105
rect 14531 17067 14716 17097
rect 14531 17063 14606 17067
rect 14531 17029 14599 17063
rect 14640 17033 14716 17067
rect 14633 17029 14716 17033
rect 14531 16995 14716 17029
rect 14531 16961 14599 16995
rect 14640 16961 14716 16995
rect 14531 16927 14716 16961
rect 14531 16893 14599 16927
rect 14633 16923 14716 16927
rect 14531 16889 14606 16893
rect 14640 16889 14716 16923
rect 14531 16859 14716 16889
rect 14531 16825 14599 16859
rect 14633 16851 14716 16859
rect 14531 16817 14606 16825
rect 14640 16817 14716 16851
rect 14531 16791 14716 16817
rect 14531 16757 14599 16791
rect 14633 16779 14716 16791
rect 14531 16745 14606 16757
rect 14640 16745 14716 16779
rect 14531 16723 14716 16745
rect 14531 16689 14599 16723
rect 14633 16707 14716 16723
rect 14531 16673 14606 16689
rect 14640 16673 14716 16707
rect 14531 16655 14716 16673
rect 14531 16621 14599 16655
rect 14633 16635 14716 16655
rect 14531 16601 14606 16621
rect 14640 16601 14716 16635
rect 14531 16587 14716 16601
rect 14531 16553 14599 16587
rect 14633 16563 14716 16587
rect 14531 16529 14606 16553
rect 14640 16529 14716 16563
rect 14531 16519 14716 16529
rect 14531 16485 14599 16519
rect 14633 16491 14716 16519
rect 14531 16457 14606 16485
rect 14640 16457 14716 16491
rect 14531 16451 14716 16457
rect 14531 16417 14599 16451
rect 14633 16419 14716 16451
rect 14531 16385 14606 16417
rect 14640 16385 14716 16419
rect 14531 16383 14716 16385
rect 14531 16349 14599 16383
rect 14633 16349 14716 16383
rect 14531 16347 14716 16349
rect 14531 16315 14606 16347
rect 14531 16281 14599 16315
rect 14640 16313 14716 16347
rect 14633 16281 14716 16313
rect 14531 16275 14716 16281
rect 14531 16247 14606 16275
rect 14531 16213 14599 16247
rect 14640 16241 14716 16275
rect 14633 16213 14716 16241
rect 14531 16203 14716 16213
rect 14531 16179 14606 16203
rect 14531 16145 14599 16179
rect 14640 16169 14716 16203
rect 14633 16145 14716 16169
rect 14531 16131 14716 16145
rect 14531 16111 14606 16131
rect 14531 16077 14599 16111
rect 14640 16097 14716 16131
rect 14633 16077 14716 16097
rect 14531 16059 14716 16077
rect 14531 16043 14606 16059
rect 14531 16009 14599 16043
rect 14640 16025 14716 16059
rect 14633 16009 14716 16025
rect 14531 15987 14716 16009
rect 14531 15975 14606 15987
rect 14531 15941 14599 15975
rect 14640 15953 14716 15987
rect 14633 15941 14716 15953
rect 14531 15915 14716 15941
rect 14531 15907 14606 15915
rect 14531 15873 14599 15907
rect 14640 15881 14716 15915
rect 14633 15873 14716 15881
rect 14531 15843 14716 15873
rect 14531 15839 14606 15843
rect 14531 15805 14599 15839
rect 14640 15809 14716 15843
rect 14633 15805 14716 15809
rect 14531 15771 14716 15805
rect 14531 15737 14599 15771
rect 14640 15737 14716 15771
rect 14531 15703 14716 15737
rect 14531 15669 14599 15703
rect 14633 15699 14716 15703
rect 14531 15665 14606 15669
rect 14640 15665 14716 15699
rect 14531 15635 14716 15665
rect 14531 15601 14599 15635
rect 14633 15627 14716 15635
rect 14531 15593 14606 15601
rect 14640 15593 14716 15627
rect 14531 15567 14716 15593
rect 14531 15533 14599 15567
rect 14633 15555 14716 15567
rect 14531 15521 14606 15533
rect 14640 15521 14716 15555
rect 14531 15499 14716 15521
rect 14531 15465 14599 15499
rect 14633 15483 14716 15499
rect 14531 15449 14606 15465
rect 14640 15449 14716 15483
rect 14531 15431 14716 15449
rect 14531 15397 14599 15431
rect 14633 15411 14716 15431
rect 14531 15377 14606 15397
rect 14640 15377 14716 15411
rect 14531 15363 14716 15377
rect 14531 15329 14599 15363
rect 14633 15339 14716 15363
rect 14531 15305 14606 15329
rect 14640 15305 14716 15339
rect 14531 15295 14716 15305
rect 14531 15261 14599 15295
rect 14633 15267 14716 15295
rect 14531 15233 14606 15261
rect 14640 15233 14716 15267
rect 14531 15227 14716 15233
rect 14531 15193 14599 15227
rect 14633 15195 14716 15227
rect 14531 15161 14606 15193
rect 14640 15161 14716 15195
rect 14531 15159 14716 15161
rect 14531 15125 14599 15159
rect 14633 15125 14716 15159
rect 14531 15123 14716 15125
rect 14531 15091 14606 15123
rect 14531 15057 14599 15091
rect 14640 15089 14716 15123
rect 14633 15057 14716 15089
rect 14531 15051 14716 15057
rect 14531 15023 14606 15051
rect 14531 14989 14599 15023
rect 14640 15017 14716 15051
rect 14633 14989 14716 15017
rect 14531 14979 14716 14989
rect 14531 14955 14606 14979
rect 14531 14921 14599 14955
rect 14640 14945 14716 14979
rect 14633 14921 14716 14945
rect 14531 14907 14716 14921
rect 14531 14887 14606 14907
rect 14531 14853 14599 14887
rect 14640 14873 14716 14907
rect 14633 14853 14716 14873
rect 14531 14835 14716 14853
rect 14531 14819 14606 14835
rect 14531 14785 14599 14819
rect 14640 14801 14716 14835
rect 14633 14785 14716 14801
rect 14531 14763 14716 14785
rect 14531 14751 14606 14763
rect 874 14723 2062 14724
rect 12874 14723 14062 14724
rect 237 14694 422 14711
rect 237 14677 312 14694
rect 237 14643 304 14677
rect 346 14660 422 14694
rect 338 14643 422 14660
rect 237 14609 422 14643
rect 237 14575 304 14609
rect 338 14575 422 14609
rect 237 14541 422 14575
rect 14531 14717 14599 14751
rect 14640 14729 14716 14763
rect 14633 14717 14716 14729
rect 14531 14691 14716 14717
rect 14531 14683 14606 14691
rect 14531 14649 14599 14683
rect 14640 14657 14716 14691
rect 14633 14649 14716 14657
rect 14531 14615 14716 14649
rect 14531 14581 14599 14615
rect 14633 14581 14716 14615
rect 14531 14541 14716 14581
rect 237 14465 14716 14541
rect 237 14431 312 14465
rect 346 14464 602 14465
rect 636 14464 2303 14465
rect 2337 14464 2375 14465
rect 2409 14464 2447 14465
rect 2481 14464 2519 14465
rect 2553 14464 2591 14465
rect 2625 14464 2663 14465
rect 2697 14464 2735 14465
rect 2769 14464 2807 14465
rect 2841 14464 2879 14465
rect 2913 14464 2951 14465
rect 2985 14464 3023 14465
rect 3057 14464 3095 14465
rect 3129 14464 3167 14465
rect 3201 14464 3239 14465
rect 3273 14464 3311 14465
rect 3345 14464 3383 14465
rect 3417 14464 3455 14465
rect 3489 14464 3527 14465
rect 3561 14464 3599 14465
rect 3633 14464 3671 14465
rect 3705 14464 3743 14465
rect 3777 14464 3815 14465
rect 3849 14464 3887 14465
rect 3921 14464 3959 14465
rect 3993 14464 4031 14465
rect 4065 14464 4103 14465
rect 4137 14464 4175 14465
rect 4209 14464 4247 14465
rect 4281 14464 4319 14465
rect 4353 14464 4391 14465
rect 4425 14464 4463 14465
rect 4497 14464 4535 14465
rect 4569 14464 4607 14465
rect 4641 14464 4679 14465
rect 4713 14464 4751 14465
rect 4785 14464 4823 14465
rect 4857 14464 4895 14465
rect 4929 14464 4967 14465
rect 5001 14464 5039 14465
rect 5073 14464 5111 14465
rect 5145 14464 5183 14465
rect 5217 14464 5255 14465
rect 5289 14464 5327 14465
rect 5361 14464 5399 14465
rect 5433 14464 5471 14465
rect 5505 14464 5543 14465
rect 5577 14464 5615 14465
rect 5649 14464 5687 14465
rect 5721 14464 5759 14465
rect 5793 14464 5831 14465
rect 5865 14464 5903 14465
rect 5937 14464 5975 14465
rect 6009 14464 6047 14465
rect 6081 14464 6119 14465
rect 6153 14464 6191 14465
rect 6225 14464 6263 14465
rect 6297 14464 6335 14465
rect 6369 14464 6407 14465
rect 6441 14464 6479 14465
rect 6513 14464 6551 14465
rect 6585 14464 6623 14465
rect 6657 14464 6695 14465
rect 6729 14464 6767 14465
rect 6801 14464 6839 14465
rect 6873 14464 6911 14465
rect 6945 14464 6983 14465
rect 7017 14464 7055 14465
rect 7089 14464 7127 14465
rect 7161 14464 7199 14465
rect 7233 14464 7271 14465
rect 7305 14464 7343 14465
rect 7377 14464 7415 14465
rect 7449 14464 7487 14465
rect 7521 14464 7559 14465
rect 7593 14464 7631 14465
rect 7665 14464 7703 14465
rect 7737 14464 7775 14465
rect 7809 14464 7847 14465
rect 7881 14464 7919 14465
rect 7953 14464 7991 14465
rect 8025 14464 8063 14465
rect 8097 14464 8135 14465
rect 8169 14464 8207 14465
rect 8241 14464 8279 14465
rect 8313 14464 8351 14465
rect 8385 14464 8423 14465
rect 8457 14464 8495 14465
rect 8529 14464 8567 14465
rect 8601 14464 8639 14465
rect 8673 14464 8711 14465
rect 8745 14464 8783 14465
rect 8817 14464 8855 14465
rect 8889 14464 8927 14465
rect 8961 14464 8999 14465
rect 9033 14464 9071 14465
rect 9105 14464 9143 14465
rect 9177 14464 9215 14465
rect 9249 14464 9287 14465
rect 9321 14464 9359 14465
rect 9393 14464 9431 14465
rect 9465 14464 9503 14465
rect 9537 14464 9575 14465
rect 9609 14464 9647 14465
rect 9681 14464 9719 14465
rect 9753 14464 9791 14465
rect 9825 14464 9863 14465
rect 9897 14464 9935 14465
rect 9969 14464 10007 14465
rect 10041 14464 10079 14465
rect 10113 14464 10151 14465
rect 10185 14464 10223 14465
rect 10257 14464 10295 14465
rect 10329 14464 10367 14465
rect 10401 14464 10439 14465
rect 10473 14464 10511 14465
rect 10545 14464 10583 14465
rect 10617 14464 10655 14465
rect 10689 14464 10727 14465
rect 10761 14464 10799 14465
rect 10833 14464 10871 14465
rect 10905 14464 10943 14465
rect 10977 14464 11015 14465
rect 11049 14464 11087 14465
rect 11121 14464 11159 14465
rect 11193 14464 11231 14465
rect 11265 14464 11303 14465
rect 11337 14464 11375 14465
rect 11409 14464 11447 14465
rect 11481 14464 11519 14465
rect 11553 14464 11591 14465
rect 11625 14464 11663 14465
rect 11697 14464 11735 14465
rect 11769 14464 11807 14465
rect 11841 14464 11879 14465
rect 11913 14464 11951 14465
rect 11985 14464 12023 14465
rect 12057 14464 12095 14465
rect 12129 14464 12167 14465
rect 12201 14464 12239 14465
rect 12273 14464 12311 14465
rect 12345 14464 12383 14465
rect 12417 14464 12455 14465
rect 12489 14464 12527 14465
rect 12561 14464 12599 14465
rect 12633 14464 14306 14465
rect 346 14431 468 14464
rect 237 14430 468 14431
rect 502 14430 536 14464
rect 570 14431 602 14464
rect 570 14430 604 14431
rect 638 14430 672 14464
rect 706 14430 740 14464
rect 774 14430 808 14464
rect 842 14430 876 14464
rect 910 14430 944 14464
rect 978 14430 1012 14464
rect 1046 14430 1080 14464
rect 1114 14430 1148 14464
rect 1182 14430 1216 14464
rect 1250 14430 1284 14464
rect 1318 14430 1352 14464
rect 1386 14430 1420 14464
rect 1454 14430 1488 14464
rect 1522 14430 1556 14464
rect 1590 14430 1624 14464
rect 1658 14430 1692 14464
rect 1726 14430 1760 14464
rect 1794 14430 1828 14464
rect 1862 14430 1896 14464
rect 1930 14430 1964 14464
rect 1998 14430 2032 14464
rect 2066 14430 2100 14464
rect 2134 14430 2168 14464
rect 2202 14430 2236 14464
rect 2270 14431 2303 14464
rect 2270 14430 2304 14431
rect 2338 14430 2372 14464
rect 2409 14431 2440 14464
rect 2481 14431 2508 14464
rect 2553 14431 2576 14464
rect 2625 14431 2644 14464
rect 2697 14431 2712 14464
rect 2769 14431 2780 14464
rect 2841 14431 2848 14464
rect 2913 14431 2916 14464
rect 2406 14430 2440 14431
rect 2474 14430 2508 14431
rect 2542 14430 2576 14431
rect 2610 14430 2644 14431
rect 2678 14430 2712 14431
rect 2746 14430 2780 14431
rect 2814 14430 2848 14431
rect 2882 14430 2916 14431
rect 2950 14431 2951 14464
rect 3018 14431 3023 14464
rect 3086 14431 3095 14464
rect 3154 14431 3167 14464
rect 3222 14431 3239 14464
rect 3290 14431 3311 14464
rect 3358 14431 3383 14464
rect 3426 14431 3455 14464
rect 3494 14431 3527 14464
rect 2950 14430 2984 14431
rect 3018 14430 3052 14431
rect 3086 14430 3120 14431
rect 3154 14430 3188 14431
rect 3222 14430 3256 14431
rect 3290 14430 3324 14431
rect 3358 14430 3392 14431
rect 3426 14430 3460 14431
rect 3494 14430 3528 14431
rect 3562 14430 3596 14464
rect 3633 14431 3664 14464
rect 3705 14431 3732 14464
rect 3777 14431 3800 14464
rect 3849 14431 3868 14464
rect 3921 14431 3936 14464
rect 3993 14431 4004 14464
rect 4065 14431 4072 14464
rect 4137 14431 4140 14464
rect 3630 14430 3664 14431
rect 3698 14430 3732 14431
rect 3766 14430 3800 14431
rect 3834 14430 3868 14431
rect 3902 14430 3936 14431
rect 3970 14430 4004 14431
rect 4038 14430 4072 14431
rect 4106 14430 4140 14431
rect 4174 14431 4175 14464
rect 4242 14431 4247 14464
rect 4310 14431 4319 14464
rect 4378 14431 4391 14464
rect 4446 14431 4463 14464
rect 4514 14431 4535 14464
rect 4582 14431 4607 14464
rect 4650 14431 4679 14464
rect 4718 14431 4751 14464
rect 4174 14430 4208 14431
rect 4242 14430 4276 14431
rect 4310 14430 4344 14431
rect 4378 14430 4412 14431
rect 4446 14430 4480 14431
rect 4514 14430 4548 14431
rect 4582 14430 4616 14431
rect 4650 14430 4684 14431
rect 4718 14430 4752 14431
rect 4786 14430 4820 14464
rect 4857 14431 4888 14464
rect 4929 14431 4956 14464
rect 5001 14431 5024 14464
rect 5073 14431 5092 14464
rect 5145 14431 5160 14464
rect 5217 14431 5228 14464
rect 5289 14431 5296 14464
rect 5361 14431 5364 14464
rect 4854 14430 4888 14431
rect 4922 14430 4956 14431
rect 4990 14430 5024 14431
rect 5058 14430 5092 14431
rect 5126 14430 5160 14431
rect 5194 14430 5228 14431
rect 5262 14430 5296 14431
rect 5330 14430 5364 14431
rect 5398 14431 5399 14464
rect 5466 14431 5471 14464
rect 5534 14431 5543 14464
rect 5602 14431 5615 14464
rect 5670 14431 5687 14464
rect 5738 14431 5759 14464
rect 5806 14431 5831 14464
rect 5874 14431 5903 14464
rect 5942 14431 5975 14464
rect 5398 14430 5432 14431
rect 5466 14430 5500 14431
rect 5534 14430 5568 14431
rect 5602 14430 5636 14431
rect 5670 14430 5704 14431
rect 5738 14430 5772 14431
rect 5806 14430 5840 14431
rect 5874 14430 5908 14431
rect 5942 14430 5976 14431
rect 6010 14430 6044 14464
rect 6081 14431 6112 14464
rect 6153 14431 6180 14464
rect 6225 14431 6248 14464
rect 6297 14431 6316 14464
rect 6369 14431 6384 14464
rect 6441 14431 6452 14464
rect 6513 14431 6520 14464
rect 6585 14431 6588 14464
rect 6078 14430 6112 14431
rect 6146 14430 6180 14431
rect 6214 14430 6248 14431
rect 6282 14430 6316 14431
rect 6350 14430 6384 14431
rect 6418 14430 6452 14431
rect 6486 14430 6520 14431
rect 6554 14430 6588 14431
rect 6622 14431 6623 14464
rect 6690 14431 6695 14464
rect 6758 14431 6767 14464
rect 6826 14431 6839 14464
rect 6894 14431 6911 14464
rect 6962 14431 6983 14464
rect 7030 14431 7055 14464
rect 7098 14431 7127 14464
rect 7166 14431 7199 14464
rect 6622 14430 6656 14431
rect 6690 14430 6724 14431
rect 6758 14430 6792 14431
rect 6826 14430 6860 14431
rect 6894 14430 6928 14431
rect 6962 14430 6996 14431
rect 7030 14430 7064 14431
rect 7098 14430 7132 14431
rect 7166 14430 7200 14431
rect 7234 14430 7268 14464
rect 7305 14431 7336 14464
rect 7377 14431 7404 14464
rect 7449 14431 7472 14464
rect 7521 14431 7540 14464
rect 7593 14431 7608 14464
rect 7665 14431 7676 14464
rect 7737 14431 7744 14464
rect 7809 14431 7812 14464
rect 7302 14430 7336 14431
rect 7370 14430 7404 14431
rect 7438 14430 7472 14431
rect 7506 14430 7540 14431
rect 7574 14430 7608 14431
rect 7642 14430 7676 14431
rect 7710 14430 7744 14431
rect 7778 14430 7812 14431
rect 7846 14431 7847 14464
rect 7914 14431 7919 14464
rect 7982 14431 7991 14464
rect 8050 14431 8063 14464
rect 8118 14431 8135 14464
rect 8186 14431 8207 14464
rect 8254 14431 8279 14464
rect 8322 14431 8351 14464
rect 8390 14431 8423 14464
rect 7846 14430 7880 14431
rect 7914 14430 7948 14431
rect 7982 14430 8016 14431
rect 8050 14430 8084 14431
rect 8118 14430 8152 14431
rect 8186 14430 8220 14431
rect 8254 14430 8288 14431
rect 8322 14430 8356 14431
rect 8390 14430 8424 14431
rect 8458 14430 8492 14464
rect 8529 14431 8560 14464
rect 8601 14431 8628 14464
rect 8673 14431 8696 14464
rect 8745 14431 8764 14464
rect 8817 14431 8832 14464
rect 8889 14431 8900 14464
rect 8961 14431 8968 14464
rect 9033 14431 9036 14464
rect 8526 14430 8560 14431
rect 8594 14430 8628 14431
rect 8662 14430 8696 14431
rect 8730 14430 8764 14431
rect 8798 14430 8832 14431
rect 8866 14430 8900 14431
rect 8934 14430 8968 14431
rect 9002 14430 9036 14431
rect 9070 14431 9071 14464
rect 9138 14431 9143 14464
rect 9206 14431 9215 14464
rect 9274 14431 9287 14464
rect 9342 14431 9359 14464
rect 9410 14431 9431 14464
rect 9478 14431 9503 14464
rect 9546 14431 9575 14464
rect 9614 14431 9647 14464
rect 9070 14430 9104 14431
rect 9138 14430 9172 14431
rect 9206 14430 9240 14431
rect 9274 14430 9308 14431
rect 9342 14430 9376 14431
rect 9410 14430 9444 14431
rect 9478 14430 9512 14431
rect 9546 14430 9580 14431
rect 9614 14430 9648 14431
rect 9682 14430 9716 14464
rect 9753 14431 9784 14464
rect 9825 14431 9852 14464
rect 9897 14431 9920 14464
rect 9969 14431 9988 14464
rect 10041 14431 10056 14464
rect 10113 14431 10124 14464
rect 10185 14431 10192 14464
rect 10257 14431 10260 14464
rect 9750 14430 9784 14431
rect 9818 14430 9852 14431
rect 9886 14430 9920 14431
rect 9954 14430 9988 14431
rect 10022 14430 10056 14431
rect 10090 14430 10124 14431
rect 10158 14430 10192 14431
rect 10226 14430 10260 14431
rect 10294 14431 10295 14464
rect 10362 14431 10367 14464
rect 10430 14431 10439 14464
rect 10498 14431 10511 14464
rect 10566 14431 10583 14464
rect 10634 14431 10655 14464
rect 10702 14431 10727 14464
rect 10770 14431 10799 14464
rect 10838 14431 10871 14464
rect 10294 14430 10328 14431
rect 10362 14430 10396 14431
rect 10430 14430 10464 14431
rect 10498 14430 10532 14431
rect 10566 14430 10600 14431
rect 10634 14430 10668 14431
rect 10702 14430 10736 14431
rect 10770 14430 10804 14431
rect 10838 14430 10872 14431
rect 10906 14430 10940 14464
rect 10977 14431 11008 14464
rect 11049 14431 11076 14464
rect 11121 14431 11144 14464
rect 11193 14431 11212 14464
rect 11265 14431 11280 14464
rect 11337 14431 11348 14464
rect 11409 14431 11416 14464
rect 11481 14431 11484 14464
rect 10974 14430 11008 14431
rect 11042 14430 11076 14431
rect 11110 14430 11144 14431
rect 11178 14430 11212 14431
rect 11246 14430 11280 14431
rect 11314 14430 11348 14431
rect 11382 14430 11416 14431
rect 11450 14430 11484 14431
rect 11518 14431 11519 14464
rect 11586 14431 11591 14464
rect 11654 14431 11663 14464
rect 11722 14431 11735 14464
rect 11790 14431 11807 14464
rect 11858 14431 11879 14464
rect 11926 14431 11951 14464
rect 11994 14431 12023 14464
rect 12062 14431 12095 14464
rect 11518 14430 11552 14431
rect 11586 14430 11620 14431
rect 11654 14430 11688 14431
rect 11722 14430 11756 14431
rect 11790 14430 11824 14431
rect 11858 14430 11892 14431
rect 11926 14430 11960 14431
rect 11994 14430 12028 14431
rect 12062 14430 12096 14431
rect 12130 14430 12164 14464
rect 12201 14431 12232 14464
rect 12273 14431 12300 14464
rect 12345 14431 12368 14464
rect 12417 14431 12436 14464
rect 12489 14431 12504 14464
rect 12561 14431 12572 14464
rect 12633 14431 12640 14464
rect 12198 14430 12232 14431
rect 12266 14430 12300 14431
rect 12334 14430 12368 14431
rect 12402 14430 12436 14431
rect 12470 14430 12504 14431
rect 12538 14430 12572 14431
rect 12606 14430 12640 14431
rect 12674 14430 12708 14464
rect 12742 14430 12776 14464
rect 12810 14430 12844 14464
rect 12878 14430 12912 14464
rect 12946 14430 12980 14464
rect 13014 14430 13048 14464
rect 13082 14430 13116 14464
rect 13150 14430 13184 14464
rect 13218 14430 13252 14464
rect 13286 14430 13320 14464
rect 13354 14430 13388 14464
rect 13422 14430 13456 14464
rect 13490 14430 13524 14464
rect 13558 14430 13592 14464
rect 13626 14430 13660 14464
rect 13694 14430 13728 14464
rect 13762 14430 13796 14464
rect 13830 14430 13864 14464
rect 13898 14430 13932 14464
rect 13966 14430 14000 14464
rect 14034 14430 14068 14464
rect 14102 14430 14136 14464
rect 14170 14430 14204 14464
rect 14238 14430 14272 14464
rect 14340 14464 14606 14465
rect 14306 14430 14340 14431
rect 14374 14430 14408 14464
rect 14442 14430 14476 14464
rect 14510 14431 14606 14464
rect 14640 14431 14716 14465
rect 14510 14430 14716 14431
rect 237 14356 14716 14430
<< viali >>
rect 312 36513 346 36547
rect 14606 36512 14640 36546
rect 548 36510 582 36511
rect 620 36510 654 36511
rect 692 36510 726 36511
rect 764 36510 798 36511
rect 836 36510 870 36511
rect 908 36510 942 36511
rect 980 36510 1014 36511
rect 1052 36510 1086 36511
rect 1124 36510 1158 36511
rect 1196 36510 1230 36511
rect 1268 36510 1302 36511
rect 1340 36510 1374 36511
rect 1412 36510 1446 36511
rect 1484 36510 1518 36511
rect 1556 36510 1590 36511
rect 1628 36510 1662 36511
rect 1700 36510 1734 36511
rect 1772 36510 1806 36511
rect 1844 36510 1878 36511
rect 1916 36510 1950 36511
rect 1988 36510 2022 36511
rect 2060 36510 2094 36511
rect 2132 36510 2166 36511
rect 2204 36510 2238 36511
rect 2276 36510 2310 36511
rect 2348 36510 2382 36511
rect 2420 36510 2454 36511
rect 2492 36510 2526 36511
rect 2564 36510 2598 36511
rect 2636 36510 2670 36511
rect 2708 36510 2742 36511
rect 2780 36510 2814 36511
rect 2852 36510 2886 36511
rect 2924 36510 2958 36511
rect 2996 36510 3030 36511
rect 3068 36510 3102 36511
rect 3140 36510 3174 36511
rect 3212 36510 3246 36511
rect 3284 36510 3318 36511
rect 3356 36510 3390 36511
rect 3428 36510 3462 36511
rect 3500 36510 3534 36511
rect 3572 36510 3606 36511
rect 3644 36510 3678 36511
rect 3716 36510 3750 36511
rect 3788 36510 3822 36511
rect 3860 36510 3894 36511
rect 3932 36510 3966 36511
rect 4004 36510 4038 36511
rect 4076 36510 4110 36511
rect 4148 36510 4182 36511
rect 4220 36510 4254 36511
rect 4292 36510 4326 36511
rect 4364 36510 4398 36511
rect 4436 36510 4470 36511
rect 4508 36510 4542 36511
rect 4580 36510 4614 36511
rect 4652 36510 4686 36511
rect 4724 36510 4758 36511
rect 4796 36510 4830 36511
rect 4868 36510 4902 36511
rect 4940 36510 4974 36511
rect 5012 36510 5046 36511
rect 5084 36510 5118 36511
rect 5156 36510 5190 36511
rect 5228 36510 5262 36511
rect 5300 36510 5334 36511
rect 5372 36510 5406 36511
rect 5444 36510 5478 36511
rect 5516 36510 5550 36511
rect 5588 36510 5622 36511
rect 5660 36510 5694 36511
rect 5732 36510 5766 36511
rect 5804 36510 5838 36511
rect 5876 36510 5910 36511
rect 5948 36510 5982 36511
rect 6020 36510 6054 36511
rect 6092 36510 6126 36511
rect 6164 36510 6198 36511
rect 6236 36510 6270 36511
rect 6308 36510 6342 36511
rect 6380 36510 6414 36511
rect 6452 36510 6486 36511
rect 6524 36510 6558 36511
rect 6596 36510 6630 36511
rect 6668 36510 6702 36511
rect 6740 36510 6774 36511
rect 6812 36510 6846 36511
rect 6884 36510 6918 36511
rect 6956 36510 6990 36511
rect 7028 36510 7062 36511
rect 7100 36510 7134 36511
rect 7172 36510 7206 36511
rect 7244 36510 7278 36511
rect 7316 36510 7350 36511
rect 7388 36510 7422 36511
rect 7460 36510 7494 36511
rect 7532 36510 7566 36511
rect 7604 36510 7638 36511
rect 7676 36510 7710 36511
rect 7748 36510 7782 36511
rect 7820 36510 7854 36511
rect 7892 36510 7926 36511
rect 7964 36510 7998 36511
rect 8036 36510 8070 36511
rect 8108 36510 8142 36511
rect 8180 36510 8214 36511
rect 8252 36510 8286 36511
rect 8324 36510 8358 36511
rect 8396 36510 8430 36511
rect 8468 36510 8502 36511
rect 8540 36510 8574 36511
rect 8612 36510 8646 36511
rect 8684 36510 8718 36511
rect 8756 36510 8790 36511
rect 8828 36510 8862 36511
rect 8900 36510 8934 36511
rect 8972 36510 9006 36511
rect 9044 36510 9078 36511
rect 9116 36510 9150 36511
rect 9188 36510 9222 36511
rect 9260 36510 9294 36511
rect 9332 36510 9366 36511
rect 9404 36510 9438 36511
rect 9476 36510 9510 36511
rect 9548 36510 9582 36511
rect 9620 36510 9654 36511
rect 9692 36510 9726 36511
rect 9764 36510 9798 36511
rect 9836 36510 9870 36511
rect 9908 36510 9942 36511
rect 9980 36510 10014 36511
rect 10052 36510 10086 36511
rect 10124 36510 10158 36511
rect 10196 36510 10230 36511
rect 10268 36510 10302 36511
rect 10340 36510 10374 36511
rect 10412 36510 10446 36511
rect 10484 36510 10518 36511
rect 10556 36510 10590 36511
rect 10628 36510 10662 36511
rect 10700 36510 10734 36511
rect 10772 36510 10806 36511
rect 10844 36510 10878 36511
rect 10916 36510 10950 36511
rect 10988 36510 11022 36511
rect 11060 36510 11094 36511
rect 11132 36510 11166 36511
rect 11204 36510 11238 36511
rect 11276 36510 11310 36511
rect 11348 36510 11382 36511
rect 11420 36510 11454 36511
rect 11492 36510 11526 36511
rect 11564 36510 11598 36511
rect 11636 36510 11670 36511
rect 11708 36510 11742 36511
rect 11780 36510 11814 36511
rect 11852 36510 11886 36511
rect 11924 36510 11958 36511
rect 11996 36510 12030 36511
rect 12068 36510 12102 36511
rect 12140 36510 12174 36511
rect 12212 36510 12246 36511
rect 12284 36510 12318 36511
rect 12356 36510 12390 36511
rect 12428 36510 12462 36511
rect 12500 36510 12534 36511
rect 12572 36510 12606 36511
rect 12644 36510 12678 36511
rect 12716 36510 12750 36511
rect 12788 36510 12822 36511
rect 12860 36510 12894 36511
rect 12932 36510 12966 36511
rect 13004 36510 13038 36511
rect 13076 36510 13110 36511
rect 13148 36510 13182 36511
rect 13220 36510 13254 36511
rect 13292 36510 13326 36511
rect 13364 36510 13398 36511
rect 13436 36510 13470 36511
rect 13508 36510 13542 36511
rect 13580 36510 13614 36511
rect 13652 36510 13686 36511
rect 13724 36510 13758 36511
rect 13796 36510 13830 36511
rect 13868 36510 13902 36511
rect 13940 36510 13974 36511
rect 14012 36510 14046 36511
rect 14084 36510 14118 36511
rect 14156 36510 14190 36511
rect 14228 36510 14262 36511
rect 14300 36510 14334 36511
rect 14372 36510 14406 36511
rect 548 36477 549 36510
rect 549 36477 582 36510
rect 620 36477 651 36510
rect 651 36477 654 36510
rect 692 36477 719 36510
rect 719 36477 726 36510
rect 764 36477 787 36510
rect 787 36477 798 36510
rect 836 36477 855 36510
rect 855 36477 870 36510
rect 908 36477 923 36510
rect 923 36477 942 36510
rect 980 36477 991 36510
rect 991 36477 1014 36510
rect 1052 36477 1059 36510
rect 1059 36477 1086 36510
rect 1124 36477 1127 36510
rect 1127 36477 1158 36510
rect 1196 36477 1229 36510
rect 1229 36477 1230 36510
rect 1268 36477 1297 36510
rect 1297 36477 1302 36510
rect 1340 36477 1365 36510
rect 1365 36477 1374 36510
rect 1412 36477 1433 36510
rect 1433 36477 1446 36510
rect 1484 36477 1501 36510
rect 1501 36477 1518 36510
rect 1556 36477 1569 36510
rect 1569 36477 1590 36510
rect 1628 36477 1637 36510
rect 1637 36477 1662 36510
rect 1700 36477 1705 36510
rect 1705 36477 1734 36510
rect 1772 36477 1773 36510
rect 1773 36477 1806 36510
rect 1844 36477 1875 36510
rect 1875 36477 1878 36510
rect 1916 36477 1943 36510
rect 1943 36477 1950 36510
rect 1988 36477 2011 36510
rect 2011 36477 2022 36510
rect 2060 36477 2079 36510
rect 2079 36477 2094 36510
rect 2132 36477 2147 36510
rect 2147 36477 2166 36510
rect 2204 36477 2215 36510
rect 2215 36477 2238 36510
rect 2276 36477 2283 36510
rect 2283 36477 2310 36510
rect 2348 36477 2351 36510
rect 2351 36477 2382 36510
rect 2420 36477 2453 36510
rect 2453 36477 2454 36510
rect 2492 36477 2521 36510
rect 2521 36477 2526 36510
rect 2564 36477 2589 36510
rect 2589 36477 2598 36510
rect 2636 36477 2657 36510
rect 2657 36477 2670 36510
rect 2708 36477 2725 36510
rect 2725 36477 2742 36510
rect 2780 36477 2793 36510
rect 2793 36477 2814 36510
rect 2852 36477 2861 36510
rect 2861 36477 2886 36510
rect 2924 36477 2929 36510
rect 2929 36477 2958 36510
rect 2996 36477 2997 36510
rect 2997 36477 3030 36510
rect 3068 36477 3099 36510
rect 3099 36477 3102 36510
rect 3140 36477 3167 36510
rect 3167 36477 3174 36510
rect 3212 36477 3235 36510
rect 3235 36477 3246 36510
rect 3284 36477 3303 36510
rect 3303 36477 3318 36510
rect 3356 36477 3371 36510
rect 3371 36477 3390 36510
rect 3428 36477 3439 36510
rect 3439 36477 3462 36510
rect 3500 36477 3507 36510
rect 3507 36477 3534 36510
rect 3572 36477 3575 36510
rect 3575 36477 3606 36510
rect 3644 36477 3677 36510
rect 3677 36477 3678 36510
rect 3716 36477 3745 36510
rect 3745 36477 3750 36510
rect 3788 36477 3813 36510
rect 3813 36477 3822 36510
rect 3860 36477 3881 36510
rect 3881 36477 3894 36510
rect 3932 36477 3949 36510
rect 3949 36477 3966 36510
rect 4004 36477 4017 36510
rect 4017 36477 4038 36510
rect 4076 36477 4085 36510
rect 4085 36477 4110 36510
rect 4148 36477 4153 36510
rect 4153 36477 4182 36510
rect 4220 36477 4221 36510
rect 4221 36477 4254 36510
rect 4292 36477 4323 36510
rect 4323 36477 4326 36510
rect 4364 36477 4391 36510
rect 4391 36477 4398 36510
rect 4436 36477 4459 36510
rect 4459 36477 4470 36510
rect 4508 36477 4527 36510
rect 4527 36477 4542 36510
rect 4580 36477 4595 36510
rect 4595 36477 4614 36510
rect 4652 36477 4663 36510
rect 4663 36477 4686 36510
rect 4724 36477 4731 36510
rect 4731 36477 4758 36510
rect 4796 36477 4799 36510
rect 4799 36477 4830 36510
rect 4868 36477 4901 36510
rect 4901 36477 4902 36510
rect 4940 36477 4969 36510
rect 4969 36477 4974 36510
rect 5012 36477 5037 36510
rect 5037 36477 5046 36510
rect 5084 36477 5105 36510
rect 5105 36477 5118 36510
rect 5156 36477 5173 36510
rect 5173 36477 5190 36510
rect 5228 36477 5241 36510
rect 5241 36477 5262 36510
rect 5300 36477 5309 36510
rect 5309 36477 5334 36510
rect 5372 36477 5377 36510
rect 5377 36477 5406 36510
rect 5444 36477 5445 36510
rect 5445 36477 5478 36510
rect 5516 36477 5547 36510
rect 5547 36477 5550 36510
rect 5588 36477 5615 36510
rect 5615 36477 5622 36510
rect 5660 36477 5683 36510
rect 5683 36477 5694 36510
rect 5732 36477 5751 36510
rect 5751 36477 5766 36510
rect 5804 36477 5819 36510
rect 5819 36477 5838 36510
rect 5876 36477 5887 36510
rect 5887 36477 5910 36510
rect 5948 36477 5955 36510
rect 5955 36477 5982 36510
rect 6020 36477 6023 36510
rect 6023 36477 6054 36510
rect 6092 36477 6125 36510
rect 6125 36477 6126 36510
rect 6164 36477 6193 36510
rect 6193 36477 6198 36510
rect 6236 36477 6261 36510
rect 6261 36477 6270 36510
rect 6308 36477 6329 36510
rect 6329 36477 6342 36510
rect 6380 36477 6397 36510
rect 6397 36477 6414 36510
rect 6452 36477 6465 36510
rect 6465 36477 6486 36510
rect 6524 36477 6533 36510
rect 6533 36477 6558 36510
rect 6596 36477 6601 36510
rect 6601 36477 6630 36510
rect 6668 36477 6669 36510
rect 6669 36477 6702 36510
rect 6740 36477 6771 36510
rect 6771 36477 6774 36510
rect 6812 36477 6839 36510
rect 6839 36477 6846 36510
rect 6884 36477 6907 36510
rect 6907 36477 6918 36510
rect 6956 36477 6975 36510
rect 6975 36477 6990 36510
rect 7028 36477 7043 36510
rect 7043 36477 7062 36510
rect 7100 36477 7111 36510
rect 7111 36477 7134 36510
rect 7172 36477 7179 36510
rect 7179 36477 7206 36510
rect 7244 36477 7247 36510
rect 7247 36477 7278 36510
rect 7316 36477 7349 36510
rect 7349 36477 7350 36510
rect 7388 36477 7417 36510
rect 7417 36477 7422 36510
rect 7460 36477 7485 36510
rect 7485 36477 7494 36510
rect 7532 36477 7553 36510
rect 7553 36477 7566 36510
rect 7604 36477 7621 36510
rect 7621 36477 7638 36510
rect 7676 36477 7689 36510
rect 7689 36477 7710 36510
rect 7748 36477 7757 36510
rect 7757 36477 7782 36510
rect 7820 36477 7825 36510
rect 7825 36477 7854 36510
rect 7892 36477 7893 36510
rect 7893 36477 7926 36510
rect 7964 36477 7995 36510
rect 7995 36477 7998 36510
rect 8036 36477 8063 36510
rect 8063 36477 8070 36510
rect 8108 36477 8131 36510
rect 8131 36477 8142 36510
rect 8180 36477 8199 36510
rect 8199 36477 8214 36510
rect 8252 36477 8267 36510
rect 8267 36477 8286 36510
rect 8324 36477 8335 36510
rect 8335 36477 8358 36510
rect 8396 36477 8403 36510
rect 8403 36477 8430 36510
rect 8468 36477 8471 36510
rect 8471 36477 8502 36510
rect 8540 36477 8573 36510
rect 8573 36477 8574 36510
rect 8612 36477 8641 36510
rect 8641 36477 8646 36510
rect 8684 36477 8709 36510
rect 8709 36477 8718 36510
rect 8756 36477 8777 36510
rect 8777 36477 8790 36510
rect 8828 36477 8845 36510
rect 8845 36477 8862 36510
rect 8900 36477 8913 36510
rect 8913 36477 8934 36510
rect 8972 36477 8981 36510
rect 8981 36477 9006 36510
rect 9044 36477 9049 36510
rect 9049 36477 9078 36510
rect 9116 36477 9117 36510
rect 9117 36477 9150 36510
rect 9188 36477 9219 36510
rect 9219 36477 9222 36510
rect 9260 36477 9287 36510
rect 9287 36477 9294 36510
rect 9332 36477 9355 36510
rect 9355 36477 9366 36510
rect 9404 36477 9423 36510
rect 9423 36477 9438 36510
rect 9476 36477 9491 36510
rect 9491 36477 9510 36510
rect 9548 36477 9559 36510
rect 9559 36477 9582 36510
rect 9620 36477 9627 36510
rect 9627 36477 9654 36510
rect 9692 36477 9695 36510
rect 9695 36477 9726 36510
rect 9764 36477 9797 36510
rect 9797 36477 9798 36510
rect 9836 36477 9865 36510
rect 9865 36477 9870 36510
rect 9908 36477 9933 36510
rect 9933 36477 9942 36510
rect 9980 36477 10001 36510
rect 10001 36477 10014 36510
rect 10052 36477 10069 36510
rect 10069 36477 10086 36510
rect 10124 36477 10137 36510
rect 10137 36477 10158 36510
rect 10196 36477 10205 36510
rect 10205 36477 10230 36510
rect 10268 36477 10273 36510
rect 10273 36477 10302 36510
rect 10340 36477 10341 36510
rect 10341 36477 10374 36510
rect 10412 36477 10443 36510
rect 10443 36477 10446 36510
rect 10484 36477 10511 36510
rect 10511 36477 10518 36510
rect 10556 36477 10579 36510
rect 10579 36477 10590 36510
rect 10628 36477 10647 36510
rect 10647 36477 10662 36510
rect 10700 36477 10715 36510
rect 10715 36477 10734 36510
rect 10772 36477 10783 36510
rect 10783 36477 10806 36510
rect 10844 36477 10851 36510
rect 10851 36477 10878 36510
rect 10916 36477 10919 36510
rect 10919 36477 10950 36510
rect 10988 36477 11021 36510
rect 11021 36477 11022 36510
rect 11060 36477 11089 36510
rect 11089 36477 11094 36510
rect 11132 36477 11157 36510
rect 11157 36477 11166 36510
rect 11204 36477 11225 36510
rect 11225 36477 11238 36510
rect 11276 36477 11293 36510
rect 11293 36477 11310 36510
rect 11348 36477 11361 36510
rect 11361 36477 11382 36510
rect 11420 36477 11429 36510
rect 11429 36477 11454 36510
rect 11492 36477 11497 36510
rect 11497 36477 11526 36510
rect 11564 36477 11565 36510
rect 11565 36477 11598 36510
rect 11636 36477 11667 36510
rect 11667 36477 11670 36510
rect 11708 36477 11735 36510
rect 11735 36477 11742 36510
rect 11780 36477 11803 36510
rect 11803 36477 11814 36510
rect 11852 36477 11871 36510
rect 11871 36477 11886 36510
rect 11924 36477 11939 36510
rect 11939 36477 11958 36510
rect 11996 36477 12007 36510
rect 12007 36477 12030 36510
rect 12068 36477 12075 36510
rect 12075 36477 12102 36510
rect 12140 36477 12143 36510
rect 12143 36477 12174 36510
rect 12212 36477 12245 36510
rect 12245 36477 12246 36510
rect 12284 36477 12313 36510
rect 12313 36477 12318 36510
rect 12356 36477 12381 36510
rect 12381 36477 12390 36510
rect 12428 36477 12449 36510
rect 12449 36477 12462 36510
rect 12500 36477 12517 36510
rect 12517 36477 12534 36510
rect 12572 36477 12585 36510
rect 12585 36477 12606 36510
rect 12644 36477 12653 36510
rect 12653 36477 12678 36510
rect 12716 36477 12721 36510
rect 12721 36477 12750 36510
rect 12788 36477 12789 36510
rect 12789 36477 12822 36510
rect 12860 36477 12891 36510
rect 12891 36477 12894 36510
rect 12932 36477 12959 36510
rect 12959 36477 12966 36510
rect 13004 36477 13027 36510
rect 13027 36477 13038 36510
rect 13076 36477 13095 36510
rect 13095 36477 13110 36510
rect 13148 36477 13163 36510
rect 13163 36477 13182 36510
rect 13220 36477 13231 36510
rect 13231 36477 13254 36510
rect 13292 36477 13299 36510
rect 13299 36477 13326 36510
rect 13364 36477 13367 36510
rect 13367 36477 13398 36510
rect 13436 36477 13469 36510
rect 13469 36477 13470 36510
rect 13508 36477 13537 36510
rect 13537 36477 13542 36510
rect 13580 36477 13605 36510
rect 13605 36477 13614 36510
rect 13652 36477 13673 36510
rect 13673 36477 13686 36510
rect 13724 36477 13741 36510
rect 13741 36477 13758 36510
rect 13796 36477 13809 36510
rect 13809 36477 13830 36510
rect 13868 36477 13877 36510
rect 13877 36477 13902 36510
rect 13940 36477 13945 36510
rect 13945 36477 13974 36510
rect 14012 36477 14013 36510
rect 14013 36477 14046 36510
rect 14084 36477 14115 36510
rect 14115 36477 14118 36510
rect 14156 36477 14183 36510
rect 14183 36477 14190 36510
rect 14228 36477 14251 36510
rect 14251 36477 14262 36510
rect 14300 36477 14319 36510
rect 14319 36477 14334 36510
rect 14372 36477 14387 36510
rect 14387 36477 14406 36510
rect 312 36441 346 36475
rect 14606 36440 14640 36474
rect 312 36267 338 36294
rect 338 36267 346 36294
rect 312 36260 346 36267
rect 312 36199 338 36222
rect 338 36199 346 36222
rect 312 36188 346 36199
rect 14606 36273 14633 36291
rect 14633 36273 14640 36291
rect 14606 36257 14640 36273
rect 312 36131 338 36150
rect 338 36131 346 36150
rect 312 36116 346 36131
rect 312 36063 338 36078
rect 338 36063 346 36078
rect 312 36044 346 36063
rect 312 35995 338 36006
rect 338 35995 346 36006
rect 312 35972 346 35995
rect 312 35927 338 35934
rect 338 35927 346 35934
rect 312 35900 346 35927
rect 312 35859 338 35862
rect 338 35859 346 35862
rect 312 35828 346 35859
rect 312 35757 346 35790
rect 312 35756 338 35757
rect 338 35756 346 35757
rect 312 35689 346 35718
rect 312 35684 338 35689
rect 338 35684 346 35689
rect 312 35621 346 35646
rect 312 35612 338 35621
rect 338 35612 346 35621
rect 312 35553 346 35574
rect 312 35540 338 35553
rect 338 35540 346 35553
rect 312 35485 346 35502
rect 312 35468 338 35485
rect 338 35468 346 35485
rect 312 35417 346 35430
rect 312 35396 338 35417
rect 338 35396 346 35417
rect 312 35349 346 35358
rect 312 35324 338 35349
rect 338 35324 346 35349
rect 312 35281 346 35286
rect 312 35252 338 35281
rect 338 35252 346 35281
rect 312 35213 346 35214
rect 312 35180 338 35213
rect 338 35180 346 35213
rect 312 35111 338 35142
rect 338 35111 346 35142
rect 312 35108 346 35111
rect 312 35043 338 35070
rect 338 35043 346 35070
rect 312 35036 346 35043
rect 312 34975 338 34998
rect 338 34975 346 34998
rect 312 34964 346 34975
rect 312 34907 338 34926
rect 338 34907 346 34926
rect 312 34892 346 34907
rect 312 34839 338 34854
rect 338 34839 346 34854
rect 312 34820 346 34839
rect 312 34771 338 34782
rect 338 34771 346 34782
rect 312 34748 346 34771
rect 312 34703 338 34710
rect 338 34703 346 34710
rect 312 34676 346 34703
rect 312 34635 338 34638
rect 338 34635 346 34638
rect 312 34604 346 34635
rect 312 34533 346 34566
rect 312 34532 338 34533
rect 338 34532 346 34533
rect 312 34465 346 34494
rect 312 34460 338 34465
rect 338 34460 346 34465
rect 312 34397 346 34422
rect 312 34388 338 34397
rect 338 34388 346 34397
rect 312 34329 346 34350
rect 312 34316 338 34329
rect 338 34316 346 34329
rect 312 34261 346 34278
rect 312 34244 338 34261
rect 338 34244 346 34261
rect 312 34193 346 34206
rect 312 34172 338 34193
rect 338 34172 346 34193
rect 312 34125 346 34134
rect 312 34100 338 34125
rect 338 34100 346 34125
rect 312 34057 346 34062
rect 312 34028 338 34057
rect 338 34028 346 34057
rect 312 33989 346 33990
rect 312 33956 338 33989
rect 338 33956 346 33989
rect 312 33887 338 33918
rect 338 33887 346 33918
rect 312 33884 346 33887
rect 312 33819 338 33846
rect 338 33819 346 33846
rect 312 33812 346 33819
rect 312 33751 338 33774
rect 338 33751 346 33774
rect 312 33740 346 33751
rect 312 33683 338 33702
rect 338 33683 346 33702
rect 312 33668 346 33683
rect 312 33615 338 33630
rect 338 33615 346 33630
rect 312 33596 346 33615
rect 312 33547 338 33558
rect 338 33547 346 33558
rect 312 33524 346 33547
rect 312 33479 338 33486
rect 338 33479 346 33486
rect 312 33452 346 33479
rect 312 33411 338 33414
rect 338 33411 346 33414
rect 312 33380 346 33411
rect 312 33309 346 33342
rect 312 33308 338 33309
rect 338 33308 346 33309
rect 312 33241 346 33270
rect 312 33236 338 33241
rect 338 33236 346 33241
rect 312 33173 346 33198
rect 312 33164 338 33173
rect 338 33164 346 33173
rect 312 33105 346 33126
rect 312 33092 338 33105
rect 338 33092 346 33105
rect 312 33037 346 33054
rect 312 33020 338 33037
rect 338 33020 346 33037
rect 312 32969 346 32982
rect 312 32948 338 32969
rect 338 32948 346 32969
rect 312 32901 346 32910
rect 312 32876 338 32901
rect 338 32876 346 32901
rect 312 32833 346 32838
rect 312 32804 338 32833
rect 338 32804 346 32833
rect 312 32765 346 32766
rect 312 32732 338 32765
rect 338 32732 346 32765
rect 312 32663 338 32694
rect 338 32663 346 32694
rect 312 32660 346 32663
rect 312 32595 338 32622
rect 338 32595 346 32622
rect 312 32588 346 32595
rect 312 32527 338 32550
rect 338 32527 346 32550
rect 312 32516 346 32527
rect 312 32459 338 32478
rect 338 32459 346 32478
rect 312 32444 346 32459
rect 312 32391 338 32406
rect 338 32391 346 32406
rect 312 32372 346 32391
rect 312 32323 338 32334
rect 338 32323 346 32334
rect 312 32300 346 32323
rect 312 32255 338 32262
rect 338 32255 346 32262
rect 312 32228 346 32255
rect 312 32187 338 32190
rect 338 32187 346 32190
rect 312 32156 346 32187
rect 312 32085 346 32118
rect 312 32084 338 32085
rect 338 32084 346 32085
rect 312 32017 346 32046
rect 312 32012 338 32017
rect 338 32012 346 32017
rect 312 31949 346 31974
rect 312 31940 338 31949
rect 338 31940 346 31949
rect 312 31881 346 31902
rect 312 31868 338 31881
rect 338 31868 346 31881
rect 312 31813 346 31830
rect 312 31796 338 31813
rect 338 31796 346 31813
rect 312 31745 346 31758
rect 312 31724 338 31745
rect 338 31724 346 31745
rect 312 31677 346 31686
rect 312 31652 338 31677
rect 338 31652 346 31677
rect 312 31609 346 31614
rect 312 31580 338 31609
rect 338 31580 346 31609
rect 312 31541 346 31542
rect 312 31508 338 31541
rect 338 31508 346 31541
rect 312 31439 338 31470
rect 338 31439 346 31470
rect 312 31436 346 31439
rect 312 31371 338 31398
rect 338 31371 346 31398
rect 312 31364 346 31371
rect 312 31303 338 31326
rect 338 31303 346 31326
rect 312 31292 346 31303
rect 312 31235 338 31254
rect 338 31235 346 31254
rect 312 31220 346 31235
rect 312 31167 338 31182
rect 338 31167 346 31182
rect 312 31148 346 31167
rect 312 31099 338 31110
rect 338 31099 346 31110
rect 312 31076 346 31099
rect 312 31031 338 31038
rect 338 31031 346 31038
rect 312 31004 346 31031
rect 312 30963 338 30966
rect 338 30963 346 30966
rect 312 30932 346 30963
rect 312 30861 346 30894
rect 312 30860 338 30861
rect 338 30860 346 30861
rect 312 30793 346 30822
rect 312 30788 338 30793
rect 338 30788 346 30793
rect 312 30725 346 30750
rect 312 30716 338 30725
rect 338 30716 346 30725
rect 312 30657 346 30678
rect 312 30644 338 30657
rect 338 30644 346 30657
rect 312 30589 346 30606
rect 312 30572 338 30589
rect 338 30572 346 30589
rect 312 30521 346 30534
rect 312 30500 338 30521
rect 338 30500 346 30521
rect 312 30453 346 30462
rect 312 30428 338 30453
rect 338 30428 346 30453
rect 312 30385 346 30390
rect 312 30356 338 30385
rect 338 30356 346 30385
rect 312 30317 346 30318
rect 312 30284 338 30317
rect 338 30284 346 30317
rect 312 30215 338 30246
rect 338 30215 346 30246
rect 312 30212 346 30215
rect 312 30147 338 30174
rect 338 30147 346 30174
rect 312 30140 346 30147
rect 312 30079 338 30102
rect 338 30079 346 30102
rect 312 30068 346 30079
rect 312 30011 338 30030
rect 338 30011 346 30030
rect 312 29996 346 30011
rect 312 29943 338 29958
rect 338 29943 346 29958
rect 312 29924 346 29943
rect 312 29875 338 29886
rect 338 29875 346 29886
rect 312 29852 346 29875
rect 312 29807 338 29814
rect 338 29807 346 29814
rect 312 29780 346 29807
rect 312 29739 338 29742
rect 338 29739 346 29742
rect 312 29708 346 29739
rect 312 29637 346 29670
rect 312 29636 338 29637
rect 338 29636 346 29637
rect 312 29569 346 29598
rect 312 29564 338 29569
rect 338 29564 346 29569
rect 312 29501 346 29526
rect 312 29492 338 29501
rect 338 29492 346 29501
rect 312 29433 346 29454
rect 312 29420 338 29433
rect 338 29420 346 29433
rect 312 29365 346 29382
rect 312 29348 338 29365
rect 338 29348 346 29365
rect 312 29297 346 29310
rect 312 29276 338 29297
rect 338 29276 346 29297
rect 312 29229 346 29238
rect 312 29204 338 29229
rect 338 29204 346 29229
rect 312 29161 346 29166
rect 312 29132 338 29161
rect 338 29132 346 29161
rect 312 29093 346 29094
rect 312 29060 338 29093
rect 338 29060 346 29093
rect 312 28991 338 29022
rect 338 28991 346 29022
rect 312 28988 346 28991
rect 312 28923 338 28950
rect 338 28923 346 28950
rect 312 28916 346 28923
rect 312 28855 338 28878
rect 338 28855 346 28878
rect 312 28844 346 28855
rect 312 28787 338 28806
rect 338 28787 346 28806
rect 312 28772 346 28787
rect 312 28719 338 28734
rect 338 28719 346 28734
rect 312 28700 346 28719
rect 312 28651 338 28662
rect 338 28651 346 28662
rect 312 28628 346 28651
rect 312 28583 338 28590
rect 338 28583 346 28590
rect 312 28556 346 28583
rect 312 28515 338 28518
rect 338 28515 346 28518
rect 312 28484 346 28515
rect 312 28413 346 28446
rect 312 28412 338 28413
rect 338 28412 346 28413
rect 312 28345 346 28374
rect 312 28340 338 28345
rect 338 28340 346 28345
rect 312 28277 346 28302
rect 312 28268 338 28277
rect 338 28268 346 28277
rect 312 28209 346 28230
rect 312 28196 338 28209
rect 338 28196 346 28209
rect 312 28141 346 28158
rect 312 28124 338 28141
rect 338 28124 346 28141
rect 312 28073 346 28086
rect 312 28052 338 28073
rect 338 28052 346 28073
rect 312 28005 346 28014
rect 312 27980 338 28005
rect 338 27980 346 28005
rect 312 27937 346 27942
rect 312 27908 338 27937
rect 338 27908 346 27937
rect 312 27869 346 27870
rect 312 27836 338 27869
rect 338 27836 346 27869
rect 312 27767 338 27798
rect 338 27767 346 27798
rect 312 27764 346 27767
rect 312 27699 338 27726
rect 338 27699 346 27726
rect 312 27692 346 27699
rect 312 27631 338 27654
rect 338 27631 346 27654
rect 312 27620 346 27631
rect 312 27563 338 27582
rect 338 27563 346 27582
rect 312 27548 346 27563
rect 312 27495 338 27510
rect 338 27495 346 27510
rect 312 27476 346 27495
rect 312 27427 338 27438
rect 338 27427 346 27438
rect 312 27404 346 27427
rect 312 27359 338 27366
rect 338 27359 346 27366
rect 312 27332 346 27359
rect 312 27291 338 27294
rect 338 27291 346 27294
rect 312 27260 346 27291
rect 312 27189 346 27222
rect 312 27188 338 27189
rect 338 27188 346 27189
rect 312 27121 346 27150
rect 312 27116 338 27121
rect 338 27116 346 27121
rect 312 27053 346 27078
rect 312 27044 338 27053
rect 338 27044 346 27053
rect 312 26985 346 27006
rect 312 26972 338 26985
rect 338 26972 346 26985
rect 312 26917 346 26934
rect 312 26900 338 26917
rect 338 26900 346 26917
rect 312 26849 346 26862
rect 312 26828 338 26849
rect 338 26828 346 26849
rect 312 26781 346 26790
rect 312 26756 338 26781
rect 338 26756 346 26781
rect 312 26713 346 26718
rect 312 26684 338 26713
rect 338 26684 346 26713
rect 312 26645 346 26646
rect 312 26612 338 26645
rect 338 26612 346 26645
rect 312 26543 338 26574
rect 338 26543 346 26574
rect 312 26540 346 26543
rect 312 26475 338 26502
rect 338 26475 346 26502
rect 312 26468 346 26475
rect 312 26407 338 26430
rect 338 26407 346 26430
rect 312 26396 346 26407
rect 312 26339 338 26358
rect 338 26339 346 26358
rect 312 26324 346 26339
rect 312 26271 338 26286
rect 338 26271 346 26286
rect 312 26252 346 26271
rect 312 26203 338 26214
rect 338 26203 346 26214
rect 312 26180 346 26203
rect 312 26135 338 26142
rect 338 26135 346 26142
rect 312 26108 346 26135
rect 312 26067 338 26070
rect 338 26067 346 26070
rect 312 26036 346 26067
rect 312 25965 346 25998
rect 312 25964 338 25965
rect 338 25964 346 25965
rect 312 25897 346 25926
rect 312 25892 338 25897
rect 338 25892 346 25897
rect 312 25829 346 25854
rect 312 25820 338 25829
rect 338 25820 346 25829
rect 312 25761 346 25782
rect 312 25748 338 25761
rect 338 25748 346 25761
rect 312 25693 346 25710
rect 312 25676 338 25693
rect 338 25676 346 25693
rect 312 25625 346 25638
rect 312 25604 338 25625
rect 338 25604 346 25625
rect 312 25557 346 25566
rect 312 25532 338 25557
rect 338 25532 346 25557
rect 312 25489 346 25494
rect 312 25460 338 25489
rect 338 25460 346 25489
rect 312 25421 346 25422
rect 312 25388 338 25421
rect 338 25388 346 25421
rect 312 25319 338 25350
rect 338 25319 346 25350
rect 312 25316 346 25319
rect 312 25251 338 25278
rect 338 25251 346 25278
rect 312 25244 346 25251
rect 312 25183 338 25206
rect 338 25183 346 25206
rect 312 25172 346 25183
rect 312 25115 338 25134
rect 338 25115 346 25134
rect 312 25100 346 25115
rect 312 25047 338 25062
rect 338 25047 346 25062
rect 312 25028 346 25047
rect 312 24979 338 24990
rect 338 24979 346 24990
rect 312 24956 346 24979
rect 312 24911 338 24918
rect 338 24911 346 24918
rect 312 24884 346 24911
rect 312 24843 338 24846
rect 338 24843 346 24846
rect 312 24812 346 24843
rect 312 24741 346 24774
rect 312 24740 338 24741
rect 338 24740 346 24741
rect 312 24673 346 24702
rect 312 24668 338 24673
rect 338 24668 346 24673
rect 312 24605 346 24630
rect 312 24596 338 24605
rect 338 24596 346 24605
rect 312 24537 346 24558
rect 312 24524 338 24537
rect 338 24524 346 24537
rect 312 24469 346 24486
rect 312 24452 338 24469
rect 338 24452 346 24469
rect 312 24401 346 24414
rect 312 24380 338 24401
rect 338 24380 346 24401
rect 312 24333 346 24342
rect 312 24308 338 24333
rect 338 24308 346 24333
rect 312 24265 346 24270
rect 312 24236 338 24265
rect 338 24236 346 24265
rect 312 24197 346 24198
rect 312 24164 338 24197
rect 338 24164 346 24197
rect 312 24095 338 24126
rect 338 24095 346 24126
rect 312 24092 346 24095
rect 312 24027 338 24054
rect 338 24027 346 24054
rect 312 24020 346 24027
rect 312 23959 338 23982
rect 338 23959 346 23982
rect 312 23948 346 23959
rect 312 23891 338 23910
rect 338 23891 346 23910
rect 312 23876 346 23891
rect 312 23823 338 23838
rect 338 23823 346 23838
rect 312 23804 346 23823
rect 312 23755 338 23766
rect 338 23755 346 23766
rect 312 23732 346 23755
rect 312 23687 338 23694
rect 338 23687 346 23694
rect 312 23660 346 23687
rect 312 23619 338 23622
rect 338 23619 346 23622
rect 312 23588 346 23619
rect 312 23517 346 23550
rect 312 23516 338 23517
rect 338 23516 346 23517
rect 312 23449 346 23478
rect 312 23444 338 23449
rect 338 23444 346 23449
rect 312 23381 346 23406
rect 312 23372 338 23381
rect 338 23372 346 23381
rect 312 23313 346 23334
rect 312 23300 338 23313
rect 338 23300 346 23313
rect 312 23245 346 23262
rect 312 23228 338 23245
rect 338 23228 346 23245
rect 312 23177 346 23190
rect 312 23156 338 23177
rect 338 23156 346 23177
rect 312 23109 346 23118
rect 312 23084 338 23109
rect 338 23084 346 23109
rect 312 23041 346 23046
rect 312 23012 338 23041
rect 338 23012 346 23041
rect 312 22973 346 22974
rect 312 22940 338 22973
rect 338 22940 346 22973
rect 312 22871 338 22902
rect 338 22871 346 22902
rect 312 22868 346 22871
rect 312 22803 338 22830
rect 338 22803 346 22830
rect 312 22796 346 22803
rect 312 22735 338 22758
rect 338 22735 346 22758
rect 312 22724 346 22735
rect 312 22667 338 22686
rect 338 22667 346 22686
rect 312 22652 346 22667
rect 312 22599 338 22614
rect 338 22599 346 22614
rect 312 22580 346 22599
rect 312 22531 338 22542
rect 338 22531 346 22542
rect 312 22508 346 22531
rect 312 22463 338 22470
rect 338 22463 346 22470
rect 312 22436 346 22463
rect 312 22395 338 22398
rect 338 22395 346 22398
rect 312 22364 346 22395
rect 312 22293 346 22326
rect 312 22292 338 22293
rect 338 22292 346 22293
rect 312 22225 346 22254
rect 312 22220 338 22225
rect 338 22220 346 22225
rect 312 22157 346 22182
rect 312 22148 338 22157
rect 338 22148 346 22157
rect 312 22089 346 22110
rect 312 22076 338 22089
rect 338 22076 346 22089
rect 312 22021 346 22038
rect 312 22004 338 22021
rect 338 22004 346 22021
rect 312 21953 346 21966
rect 312 21932 338 21953
rect 338 21932 346 21953
rect 312 21885 346 21894
rect 312 21860 338 21885
rect 338 21860 346 21885
rect 312 21817 346 21822
rect 312 21788 338 21817
rect 338 21788 346 21817
rect 312 21749 346 21750
rect 312 21716 338 21749
rect 338 21716 346 21749
rect 312 21647 338 21678
rect 338 21647 346 21678
rect 312 21644 346 21647
rect 312 21579 338 21606
rect 338 21579 346 21606
rect 312 21572 346 21579
rect 312 21511 338 21534
rect 338 21511 346 21534
rect 312 21500 346 21511
rect 312 21443 338 21462
rect 338 21443 346 21462
rect 312 21428 346 21443
rect 312 21375 338 21390
rect 338 21375 346 21390
rect 312 21356 346 21375
rect 312 21307 338 21318
rect 338 21307 346 21318
rect 312 21284 346 21307
rect 312 21239 338 21246
rect 338 21239 346 21246
rect 312 21212 346 21239
rect 312 21171 338 21174
rect 338 21171 346 21174
rect 312 21140 346 21171
rect 312 21069 346 21102
rect 312 21068 338 21069
rect 338 21068 346 21069
rect 312 21001 346 21030
rect 312 20996 338 21001
rect 338 20996 346 21001
rect 312 20933 346 20958
rect 312 20924 338 20933
rect 338 20924 346 20933
rect 312 20865 346 20886
rect 312 20852 338 20865
rect 338 20852 346 20865
rect 312 20797 346 20814
rect 312 20780 338 20797
rect 338 20780 346 20797
rect 312 20729 346 20742
rect 312 20708 338 20729
rect 338 20708 346 20729
rect 312 20661 346 20670
rect 312 20636 338 20661
rect 338 20636 346 20661
rect 312 20593 346 20598
rect 312 20564 338 20593
rect 338 20564 346 20593
rect 312 20525 346 20526
rect 312 20492 338 20525
rect 338 20492 346 20525
rect 312 20423 338 20454
rect 338 20423 346 20454
rect 312 20420 346 20423
rect 312 20355 338 20382
rect 338 20355 346 20382
rect 312 20348 346 20355
rect 312 20287 338 20310
rect 338 20287 346 20310
rect 312 20276 346 20287
rect 312 20219 338 20238
rect 338 20219 346 20238
rect 312 20204 346 20219
rect 312 20151 338 20166
rect 338 20151 346 20166
rect 312 20132 346 20151
rect 312 20083 338 20094
rect 338 20083 346 20094
rect 312 20060 346 20083
rect 312 20015 338 20022
rect 338 20015 346 20022
rect 312 19988 346 20015
rect 312 19947 338 19950
rect 338 19947 346 19950
rect 312 19916 346 19947
rect 312 19845 346 19878
rect 312 19844 338 19845
rect 338 19844 346 19845
rect 312 19777 346 19806
rect 312 19772 338 19777
rect 338 19772 346 19777
rect 312 19709 346 19734
rect 312 19700 338 19709
rect 338 19700 346 19709
rect 312 19641 346 19662
rect 312 19628 338 19641
rect 338 19628 346 19641
rect 312 19573 346 19590
rect 312 19556 338 19573
rect 338 19556 346 19573
rect 312 19505 346 19518
rect 312 19484 338 19505
rect 338 19484 346 19505
rect 312 19437 346 19446
rect 312 19412 338 19437
rect 338 19412 346 19437
rect 312 19369 346 19374
rect 312 19340 338 19369
rect 338 19340 346 19369
rect 312 19301 346 19302
rect 312 19268 338 19301
rect 338 19268 346 19301
rect 312 19199 338 19230
rect 338 19199 346 19230
rect 312 19196 346 19199
rect 312 19131 338 19158
rect 338 19131 346 19158
rect 312 19124 346 19131
rect 312 19063 338 19086
rect 338 19063 346 19086
rect 312 19052 346 19063
rect 312 18995 338 19014
rect 338 18995 346 19014
rect 312 18980 346 18995
rect 312 18927 338 18942
rect 338 18927 346 18942
rect 312 18908 346 18927
rect 312 18859 338 18870
rect 338 18859 346 18870
rect 312 18836 346 18859
rect 312 18791 338 18798
rect 338 18791 346 18798
rect 312 18764 346 18791
rect 312 18723 338 18726
rect 338 18723 346 18726
rect 312 18692 346 18723
rect 312 18621 346 18654
rect 312 18620 338 18621
rect 338 18620 346 18621
rect 312 18553 346 18582
rect 312 18548 338 18553
rect 338 18548 346 18553
rect 312 18485 346 18510
rect 312 18476 338 18485
rect 338 18476 346 18485
rect 312 18417 346 18438
rect 312 18404 338 18417
rect 338 18404 346 18417
rect 312 18349 346 18366
rect 312 18332 338 18349
rect 338 18332 346 18349
rect 312 18281 346 18294
rect 312 18260 338 18281
rect 338 18260 346 18281
rect 312 18213 346 18222
rect 312 18188 338 18213
rect 338 18188 346 18213
rect 312 18145 346 18150
rect 312 18116 338 18145
rect 338 18116 346 18145
rect 312 18077 346 18078
rect 312 18044 338 18077
rect 338 18044 346 18077
rect 312 17975 338 18006
rect 338 17975 346 18006
rect 312 17972 346 17975
rect 312 17907 338 17934
rect 338 17907 346 17934
rect 312 17900 346 17907
rect 312 17839 338 17862
rect 338 17839 346 17862
rect 312 17828 346 17839
rect 312 17771 338 17790
rect 338 17771 346 17790
rect 312 17756 346 17771
rect 312 17703 338 17718
rect 338 17703 346 17718
rect 312 17684 346 17703
rect 312 17635 338 17646
rect 338 17635 346 17646
rect 312 17612 346 17635
rect 312 17567 338 17574
rect 338 17567 346 17574
rect 312 17540 346 17567
rect 312 17499 338 17502
rect 338 17499 346 17502
rect 312 17468 346 17499
rect 312 17397 346 17430
rect 312 17396 338 17397
rect 338 17396 346 17397
rect 312 17329 346 17358
rect 312 17324 338 17329
rect 338 17324 346 17329
rect 312 17261 346 17286
rect 312 17252 338 17261
rect 338 17252 346 17261
rect 312 17193 346 17214
rect 312 17180 338 17193
rect 338 17180 346 17193
rect 312 17125 346 17142
rect 312 17108 338 17125
rect 338 17108 346 17125
rect 312 17057 346 17070
rect 312 17036 338 17057
rect 338 17036 346 17057
rect 312 16989 346 16998
rect 312 16964 338 16989
rect 338 16964 346 16989
rect 312 16921 346 16926
rect 312 16892 338 16921
rect 338 16892 346 16921
rect 312 16853 346 16854
rect 312 16820 338 16853
rect 338 16820 346 16853
rect 312 16751 338 16782
rect 338 16751 346 16782
rect 312 16748 346 16751
rect 312 16683 338 16710
rect 338 16683 346 16710
rect 312 16676 346 16683
rect 312 16615 338 16638
rect 338 16615 346 16638
rect 312 16604 346 16615
rect 312 16547 338 16566
rect 338 16547 346 16566
rect 312 16532 346 16547
rect 312 16479 338 16494
rect 338 16479 346 16494
rect 312 16460 346 16479
rect 312 16411 338 16422
rect 338 16411 346 16422
rect 312 16388 346 16411
rect 312 16343 338 16350
rect 338 16343 346 16350
rect 312 16316 346 16343
rect 312 16275 338 16278
rect 338 16275 346 16278
rect 312 16244 346 16275
rect 312 16173 346 16206
rect 312 16172 338 16173
rect 338 16172 346 16173
rect 312 16105 346 16134
rect 312 16100 338 16105
rect 338 16100 346 16105
rect 312 16037 346 16062
rect 312 16028 338 16037
rect 338 16028 346 16037
rect 312 15969 346 15990
rect 312 15956 338 15969
rect 338 15956 346 15969
rect 312 15901 346 15918
rect 312 15884 338 15901
rect 338 15884 346 15901
rect 312 15833 346 15846
rect 312 15812 338 15833
rect 338 15812 346 15833
rect 312 15765 346 15774
rect 312 15740 338 15765
rect 338 15740 346 15765
rect 312 15697 346 15702
rect 312 15668 338 15697
rect 338 15668 346 15697
rect 312 15629 346 15630
rect 312 15596 338 15629
rect 338 15596 346 15629
rect 312 15527 338 15558
rect 338 15527 346 15558
rect 312 15524 346 15527
rect 312 15459 338 15486
rect 338 15459 346 15486
rect 312 15452 346 15459
rect 312 15391 338 15414
rect 338 15391 346 15414
rect 312 15380 346 15391
rect 312 15323 338 15342
rect 338 15323 346 15342
rect 312 15308 346 15323
rect 312 15255 338 15270
rect 338 15255 346 15270
rect 312 15236 346 15255
rect 312 15187 338 15198
rect 338 15187 346 15198
rect 312 15164 346 15187
rect 312 15119 338 15126
rect 338 15119 346 15126
rect 312 15092 346 15119
rect 312 15051 338 15054
rect 338 15051 346 15054
rect 312 15020 346 15051
rect 312 14949 346 14982
rect 312 14948 338 14949
rect 338 14948 346 14949
rect 312 14881 346 14910
rect 312 14876 338 14881
rect 338 14876 346 14881
rect 312 14813 346 14838
rect 312 14804 338 14813
rect 338 14804 346 14813
rect 312 14745 346 14766
rect 312 14732 338 14745
rect 338 14732 346 14745
rect 1001 35982 1035 36016
rect 1073 35982 1107 36016
rect 1145 35982 1179 36016
rect 1217 35982 1251 36016
rect 1289 35982 1323 36016
rect 1361 35982 1395 36016
rect 1433 35982 1467 36016
rect 1505 35982 1539 36016
rect 1577 35982 1611 36016
rect 1649 35982 1683 36016
rect 1721 35982 1755 36016
rect 1793 35982 1827 36016
rect 1865 35982 1899 36016
rect 1937 35982 1971 36016
rect 2009 35982 2043 36016
rect 2081 35982 2115 36016
rect 2153 35982 2187 36016
rect 2225 35982 2259 36016
rect 2297 35982 2331 36016
rect 2369 35982 2403 36016
rect 2441 35982 2475 36016
rect 2513 35982 2547 36016
rect 2585 35982 2619 36016
rect 2657 35982 2691 36016
rect 2729 35982 2763 36016
rect 2801 35982 2835 36016
rect 2873 35982 2907 36016
rect 2945 35982 2979 36016
rect 3017 35982 3051 36016
rect 3089 35982 3123 36016
rect 3161 35982 3195 36016
rect 3233 35982 3267 36016
rect 3305 35982 3339 36016
rect 3377 35982 3411 36016
rect 3449 35982 3483 36016
rect 3521 35982 3555 36016
rect 3593 35982 3627 36016
rect 3665 35982 3699 36016
rect 3737 35982 3771 36016
rect 3809 35982 3843 36016
rect 3881 35982 3915 36016
rect 3953 35982 3987 36016
rect 4025 35982 4059 36016
rect 4097 35982 4131 36016
rect 4169 35982 4203 36016
rect 4241 35982 4275 36016
rect 4313 35982 4347 36016
rect 4385 35982 4419 36016
rect 4457 35982 4491 36016
rect 4529 35982 4563 36016
rect 4601 35982 4635 36016
rect 4673 35982 4707 36016
rect 4745 35982 4779 36016
rect 4817 35982 4851 36016
rect 4889 35982 4923 36016
rect 4961 35982 4995 36016
rect 5033 35982 5067 36016
rect 5105 35982 5139 36016
rect 5177 35982 5211 36016
rect 5249 35982 5283 36016
rect 5321 35982 5355 36016
rect 5393 35982 5427 36016
rect 5465 35982 5499 36016
rect 5537 35982 5571 36016
rect 5609 35982 5643 36016
rect 5681 35982 5715 36016
rect 5753 35982 5787 36016
rect 5825 35982 5859 36016
rect 5897 35982 5931 36016
rect 5969 35982 6003 36016
rect 6041 35982 6075 36016
rect 6113 35982 6147 36016
rect 6185 35982 6219 36016
rect 6257 35982 6291 36016
rect 6329 35982 6363 36016
rect 6401 35982 6435 36016
rect 6473 35982 6507 36016
rect 6545 35982 6579 36016
rect 6617 35982 6651 36016
rect 6689 35982 6723 36016
rect 6761 35982 6795 36016
rect 6833 35982 6867 36016
rect 6905 35982 6939 36016
rect 6977 35982 7011 36016
rect 7049 35982 7083 36016
rect 7121 35982 7155 36016
rect 7193 35982 7227 36016
rect 7265 35982 7299 36016
rect 7337 35982 7371 36016
rect 7409 35982 7443 36016
rect 7481 35982 7515 36016
rect 7553 35982 7587 36016
rect 7625 35982 7659 36016
rect 7697 35982 7731 36016
rect 7769 35982 7803 36016
rect 7841 35982 7875 36016
rect 7913 35982 7947 36016
rect 7985 35982 8019 36016
rect 8057 35982 8091 36016
rect 8129 35982 8163 36016
rect 8201 35982 8235 36016
rect 8273 35982 8307 36016
rect 8345 35982 8379 36016
rect 8417 35982 8451 36016
rect 8489 35982 8523 36016
rect 8561 35982 8595 36016
rect 8633 35982 8667 36016
rect 8705 35982 8739 36016
rect 8777 35982 8811 36016
rect 8849 35982 8883 36016
rect 8921 35982 8955 36016
rect 8993 35982 9027 36016
rect 9065 35982 9099 36016
rect 9137 35982 9171 36016
rect 9209 35982 9243 36016
rect 9281 35982 9315 36016
rect 9353 35982 9387 36016
rect 9425 35982 9459 36016
rect 9497 35982 9531 36016
rect 9569 35982 9603 36016
rect 9641 35982 9675 36016
rect 9713 35982 9747 36016
rect 9785 35982 9819 36016
rect 9857 35982 9891 36016
rect 9929 35982 9963 36016
rect 10001 35982 10035 36016
rect 10073 35982 10107 36016
rect 10145 35982 10179 36016
rect 10217 35982 10251 36016
rect 10289 35982 10323 36016
rect 10361 35982 10395 36016
rect 10433 35982 10467 36016
rect 10505 35982 10539 36016
rect 10577 35982 10611 36016
rect 10649 35982 10683 36016
rect 10721 35982 10755 36016
rect 10793 35982 10827 36016
rect 10865 35982 10899 36016
rect 10937 35982 10971 36016
rect 11009 35982 11043 36016
rect 11081 35982 11115 36016
rect 11153 35982 11187 36016
rect 11225 35982 11259 36016
rect 11297 35982 11331 36016
rect 11369 35982 11403 36016
rect 11441 35982 11475 36016
rect 11513 35982 11547 36016
rect 11585 35982 11619 36016
rect 11657 35982 11691 36016
rect 11729 35982 11763 36016
rect 11801 35982 11835 36016
rect 11873 35982 11907 36016
rect 11945 35982 11979 36016
rect 12017 35982 12051 36016
rect 12089 35982 12123 36016
rect 12161 35982 12195 36016
rect 12233 35982 12267 36016
rect 12305 35982 12339 36016
rect 12377 35982 12411 36016
rect 12449 35982 12483 36016
rect 12521 35982 12555 36016
rect 12593 35982 12627 36016
rect 12665 35982 12699 36016
rect 12737 35982 12771 36016
rect 12809 35982 12843 36016
rect 12881 35982 12915 36016
rect 12953 35982 12987 36016
rect 13025 35982 13059 36016
rect 13097 35982 13131 36016
rect 13169 35982 13203 36016
rect 13241 35982 13275 36016
rect 13313 35982 13347 36016
rect 13385 35982 13419 36016
rect 13457 35982 13491 36016
rect 13529 35982 13563 36016
rect 13601 35982 13635 36016
rect 13673 35982 13707 36016
rect 13745 35982 13779 36016
rect 13817 35982 13851 36016
rect 13889 35982 13923 36016
rect 13961 35982 13995 36016
rect 799 35879 833 35913
rect 799 35807 833 35841
rect 14114 35800 14148 35834
rect 799 35735 833 35769
rect 14114 35728 14148 35762
rect 799 35663 833 35697
rect 14114 35656 14148 35690
rect 799 35591 833 35625
rect 14114 35584 14148 35618
rect 799 35519 833 35553
rect 14114 35512 14148 35546
rect 799 35447 833 35481
rect 14114 35440 14148 35474
rect 799 35375 833 35409
rect 14114 35368 14148 35402
rect 799 35303 833 35337
rect 14114 35296 14148 35330
rect 799 35231 833 35265
rect 14114 35224 14148 35258
rect 799 35159 833 35193
rect 14114 35152 14148 35186
rect 799 35087 833 35121
rect 14114 35080 14148 35114
rect 799 35015 833 35049
rect 14114 35008 14148 35042
rect 799 34943 833 34977
rect 14114 34936 14148 34970
rect 799 34871 833 34905
rect 14114 34864 14148 34898
rect 799 34799 833 34833
rect 799 34727 833 34761
rect 14114 34792 14148 34826
rect 799 34655 833 34689
rect 799 34583 833 34617
rect 799 34511 833 34545
rect 799 34439 833 34473
rect 799 34367 833 34401
rect 799 34295 833 34329
rect 799 34223 833 34257
rect 799 34151 833 34185
rect 799 34079 833 34113
rect 799 34007 833 34041
rect 799 33935 833 33969
rect 799 33863 833 33897
rect 799 33791 833 33825
rect 799 33719 833 33753
rect 799 33647 833 33681
rect 799 33575 833 33609
rect 799 33503 833 33537
rect 799 33431 833 33465
rect 799 33359 833 33393
rect 799 33287 833 33321
rect 799 33215 833 33249
rect 799 33143 833 33177
rect 799 33071 833 33105
rect 799 32999 833 33033
rect 799 32927 833 32961
rect 799 32855 833 32889
rect 799 32783 833 32817
rect 799 32711 833 32745
rect 799 32639 833 32673
rect 799 32567 833 32601
rect 799 32495 833 32529
rect 799 32423 833 32457
rect 799 32351 833 32385
rect 799 32279 833 32313
rect 799 32207 833 32241
rect 799 32135 833 32169
rect 799 32063 833 32097
rect 799 31991 833 32025
rect 799 31919 833 31953
rect 799 31847 833 31881
rect 799 31775 833 31809
rect 799 31703 833 31737
rect 799 31631 833 31665
rect 799 31559 833 31593
rect 799 31487 833 31521
rect 799 31415 833 31449
rect 799 31343 833 31377
rect 799 31271 833 31305
rect 799 31199 833 31233
rect 799 31127 833 31161
rect 799 31055 833 31089
rect 799 30983 833 31017
rect 799 30911 833 30945
rect 799 30839 833 30873
rect 799 30767 833 30801
rect 799 30695 833 30729
rect 799 30623 833 30657
rect 799 30551 833 30585
rect 799 30479 833 30513
rect 799 30407 833 30441
rect 799 30335 833 30369
rect 799 30263 833 30297
rect 799 30191 833 30225
rect 799 30119 833 30153
rect 799 30047 833 30081
rect 799 29975 833 30009
rect 799 29903 833 29937
rect 799 29831 833 29865
rect 799 29759 833 29793
rect 799 29687 833 29721
rect 799 29615 833 29649
rect 799 29543 833 29577
rect 799 29471 833 29505
rect 799 29399 833 29433
rect 799 29327 833 29361
rect 799 29255 833 29289
rect 799 29183 833 29217
rect 799 29111 833 29145
rect 799 29039 833 29073
rect 799 28967 833 29001
rect 799 28895 833 28929
rect 799 28823 833 28857
rect 799 28751 833 28785
rect 799 28679 833 28713
rect 799 28607 833 28641
rect 799 28535 833 28569
rect 799 28463 833 28497
rect 799 28391 833 28425
rect 799 28319 833 28353
rect 799 28247 833 28281
rect 799 28175 833 28209
rect 799 28103 833 28137
rect 799 28031 833 28065
rect 799 27959 833 27993
rect 799 27887 833 27921
rect 799 27815 833 27849
rect 799 27743 833 27777
rect 799 27671 833 27705
rect 799 27599 833 27633
rect 799 27527 833 27561
rect 799 27455 833 27489
rect 799 27383 833 27417
rect 799 27311 833 27345
rect 799 27239 833 27273
rect 799 27167 833 27201
rect 799 27095 833 27129
rect 799 27023 833 27057
rect 799 26951 833 26985
rect 799 26879 833 26913
rect 799 26807 833 26841
rect 799 26735 833 26769
rect 799 26663 833 26697
rect 799 26591 833 26625
rect 799 26519 833 26553
rect 799 26447 833 26481
rect 799 26375 833 26409
rect 799 26303 833 26337
rect 799 26231 833 26265
rect 799 26159 833 26193
rect 799 26087 833 26121
rect 799 26015 833 26049
rect 799 25943 833 25977
rect 799 25871 833 25905
rect 799 25799 833 25833
rect 799 25727 833 25761
rect 799 25655 833 25689
rect 799 25583 833 25617
rect 799 25511 833 25545
rect 799 25439 833 25473
rect 799 25367 833 25401
rect 799 25295 833 25329
rect 799 25223 833 25257
rect 799 25151 833 25185
rect 799 25079 833 25113
rect 799 25007 833 25041
rect 799 24935 833 24969
rect 799 24863 833 24897
rect 799 24791 833 24825
rect 799 24719 833 24753
rect 799 24647 833 24681
rect 799 24575 833 24609
rect 799 24503 833 24537
rect 799 24431 833 24465
rect 799 24359 833 24393
rect 799 24287 833 24321
rect 799 24215 833 24249
rect 799 24143 833 24177
rect 799 24071 833 24105
rect 799 23999 833 24033
rect 799 23927 833 23961
rect 799 23855 833 23889
rect 799 23783 833 23817
rect 799 23711 833 23745
rect 799 23639 833 23673
rect 799 23567 833 23601
rect 799 23495 833 23529
rect 799 23423 833 23457
rect 799 23351 833 23385
rect 799 23279 833 23313
rect 799 23207 833 23241
rect 799 23135 833 23169
rect 799 23063 833 23097
rect 799 22991 833 23025
rect 799 22919 833 22953
rect 799 22847 833 22881
rect 799 22775 833 22809
rect 799 22703 833 22737
rect 799 22631 833 22665
rect 799 22559 833 22593
rect 799 22487 833 22521
rect 799 22415 833 22449
rect 799 22343 833 22377
rect 799 22271 833 22305
rect 799 22199 833 22233
rect 799 22127 833 22161
rect 799 22055 833 22089
rect 799 21983 833 22017
rect 799 21911 833 21945
rect 799 21839 833 21873
rect 799 21767 833 21801
rect 799 21695 833 21729
rect 799 21623 833 21657
rect 799 21551 833 21585
rect 799 21479 833 21513
rect 799 21407 833 21441
rect 799 21335 833 21369
rect 799 21263 833 21297
rect 799 21191 833 21225
rect 799 21119 833 21153
rect 799 21047 833 21081
rect 799 20975 833 21009
rect 799 20903 833 20937
rect 799 20831 833 20865
rect 799 20759 833 20793
rect 799 20687 833 20721
rect 799 20615 833 20649
rect 799 20543 833 20577
rect 799 20471 833 20505
rect 799 20399 833 20433
rect 799 20327 833 20361
rect 799 20255 833 20289
rect 799 20183 833 20217
rect 799 20111 833 20145
rect 799 20039 833 20073
rect 799 19967 833 20001
rect 799 19895 833 19929
rect 799 19823 833 19857
rect 799 19751 833 19785
rect 799 19679 833 19713
rect 799 19607 833 19641
rect 799 19535 833 19569
rect 799 19463 833 19497
rect 799 19391 833 19425
rect 799 19319 833 19353
rect 799 19247 833 19281
rect 799 19175 833 19209
rect 799 19103 833 19137
rect 799 19031 833 19065
rect 799 18959 833 18993
rect 799 18887 833 18921
rect 799 18815 833 18849
rect 799 18743 833 18777
rect 799 18671 833 18705
rect 799 18599 833 18633
rect 799 18527 833 18561
rect 799 18455 833 18489
rect 799 18383 833 18417
rect 799 18311 833 18345
rect 799 18239 833 18273
rect 799 18167 833 18201
rect 799 18095 833 18129
rect 799 18023 833 18057
rect 799 17951 833 17985
rect 799 17879 833 17913
rect 799 17807 833 17841
rect 799 17735 833 17769
rect 799 17663 833 17697
rect 799 17591 833 17625
rect 799 17519 833 17553
rect 799 17447 833 17481
rect 799 17375 833 17409
rect 799 17303 833 17337
rect 799 17231 833 17265
rect 799 17159 833 17193
rect 799 17087 833 17121
rect 799 17015 833 17049
rect 799 16943 833 16977
rect 799 16871 833 16905
rect 799 16799 833 16833
rect 799 16727 833 16761
rect 799 16655 833 16689
rect 799 16583 833 16617
rect 799 16511 833 16545
rect 799 16439 833 16473
rect 799 16367 833 16401
rect 799 16295 833 16329
rect 799 16223 833 16257
rect 799 16151 833 16185
rect 799 16079 833 16113
rect 799 16007 833 16041
rect 799 15935 833 15969
rect 799 15863 833 15897
rect 799 15791 833 15825
rect 799 15719 833 15753
rect 799 15647 833 15681
rect 799 15575 833 15609
rect 799 15503 833 15537
rect 799 15431 833 15465
rect 799 15359 833 15393
rect 799 15287 833 15321
rect 799 15215 833 15249
rect 1293 34658 1297 34692
rect 1297 34658 1327 34692
rect 1365 34658 1399 34692
rect 1437 34658 1467 34692
rect 1467 34658 1471 34692
rect 1509 34658 1535 34692
rect 1535 34658 1543 34692
rect 1581 34658 1603 34692
rect 1603 34658 1615 34692
rect 1653 34658 1671 34692
rect 1671 34658 1687 34692
rect 1725 34658 1739 34692
rect 1739 34658 1759 34692
rect 1797 34658 1807 34692
rect 1807 34658 1831 34692
rect 1869 34658 1875 34692
rect 1875 34658 1903 34692
rect 1941 34658 1943 34692
rect 1943 34658 1975 34692
rect 2013 34658 2045 34692
rect 2045 34658 2047 34692
rect 2085 34658 2113 34692
rect 2113 34658 2119 34692
rect 2157 34658 2181 34692
rect 2181 34658 2191 34692
rect 2229 34658 2249 34692
rect 2249 34658 2263 34692
rect 2301 34658 2317 34692
rect 2317 34658 2335 34692
rect 2373 34658 2385 34692
rect 2385 34658 2407 34692
rect 2445 34658 2453 34692
rect 2453 34658 2479 34692
rect 2517 34658 2521 34692
rect 2521 34658 2551 34692
rect 2589 34658 2623 34692
rect 2661 34658 2691 34692
rect 2691 34658 2695 34692
rect 2733 34658 2759 34692
rect 2759 34658 2767 34692
rect 2805 34658 2827 34692
rect 2827 34658 2839 34692
rect 2877 34658 2895 34692
rect 2895 34658 2911 34692
rect 2949 34658 2963 34692
rect 2963 34658 2983 34692
rect 3021 34658 3031 34692
rect 3031 34658 3055 34692
rect 3093 34658 3099 34692
rect 3099 34658 3127 34692
rect 3165 34658 3167 34692
rect 3167 34658 3199 34692
rect 3237 34658 3269 34692
rect 3269 34658 3271 34692
rect 3309 34658 3337 34692
rect 3337 34658 3343 34692
rect 3381 34658 3405 34692
rect 3405 34658 3415 34692
rect 3453 34658 3473 34692
rect 3473 34658 3487 34692
rect 3525 34658 3541 34692
rect 3541 34658 3559 34692
rect 3597 34658 3609 34692
rect 3609 34658 3631 34692
rect 3669 34658 3677 34692
rect 3677 34658 3703 34692
rect 3741 34658 3745 34692
rect 3745 34658 3775 34692
rect 3813 34658 3847 34692
rect 3885 34658 3915 34692
rect 3915 34658 3919 34692
rect 3957 34658 3983 34692
rect 3983 34658 3991 34692
rect 4029 34658 4051 34692
rect 4051 34658 4063 34692
rect 4101 34658 4119 34692
rect 4119 34658 4135 34692
rect 4173 34658 4187 34692
rect 4187 34658 4207 34692
rect 4245 34658 4255 34692
rect 4255 34658 4279 34692
rect 4317 34658 4323 34692
rect 4323 34658 4351 34692
rect 4389 34658 4391 34692
rect 4391 34658 4423 34692
rect 4461 34658 4493 34692
rect 4493 34658 4495 34692
rect 4533 34658 4561 34692
rect 4561 34658 4567 34692
rect 4605 34658 4629 34692
rect 4629 34658 4639 34692
rect 4677 34658 4697 34692
rect 4697 34658 4711 34692
rect 4749 34658 4765 34692
rect 4765 34658 4783 34692
rect 4821 34658 4833 34692
rect 4833 34658 4855 34692
rect 4893 34658 4901 34692
rect 4901 34658 4927 34692
rect 4965 34658 4969 34692
rect 4969 34658 4999 34692
rect 5037 34658 5071 34692
rect 5109 34658 5139 34692
rect 5139 34658 5143 34692
rect 5181 34658 5207 34692
rect 5207 34658 5215 34692
rect 5253 34658 5275 34692
rect 5275 34658 5287 34692
rect 5325 34658 5343 34692
rect 5343 34658 5359 34692
rect 5397 34658 5411 34692
rect 5411 34658 5431 34692
rect 5469 34658 5479 34692
rect 5479 34658 5503 34692
rect 5541 34658 5547 34692
rect 5547 34658 5575 34692
rect 5613 34658 5615 34692
rect 5615 34658 5647 34692
rect 5685 34658 5717 34692
rect 5717 34658 5719 34692
rect 5757 34658 5785 34692
rect 5785 34658 5791 34692
rect 5829 34658 5853 34692
rect 5853 34658 5863 34692
rect 5901 34658 5921 34692
rect 5921 34658 5935 34692
rect 5973 34658 5989 34692
rect 5989 34658 6007 34692
rect 6045 34658 6057 34692
rect 6057 34658 6079 34692
rect 6117 34658 6125 34692
rect 6125 34658 6151 34692
rect 6189 34658 6193 34692
rect 6193 34658 6223 34692
rect 6261 34658 6295 34692
rect 6333 34658 6363 34692
rect 6363 34658 6367 34692
rect 6405 34658 6431 34692
rect 6431 34658 6439 34692
rect 6477 34658 6499 34692
rect 6499 34658 6511 34692
rect 6549 34658 6567 34692
rect 6567 34658 6583 34692
rect 6621 34658 6635 34692
rect 6635 34658 6655 34692
rect 6693 34658 6703 34692
rect 6703 34658 6727 34692
rect 6765 34658 6771 34692
rect 6771 34658 6799 34692
rect 6837 34658 6839 34692
rect 6839 34658 6871 34692
rect 6909 34658 6941 34692
rect 6941 34658 6943 34692
rect 6981 34658 7009 34692
rect 7009 34658 7015 34692
rect 7053 34658 7077 34692
rect 7077 34658 7087 34692
rect 7125 34658 7145 34692
rect 7145 34658 7159 34692
rect 7197 34658 7213 34692
rect 7213 34658 7231 34692
rect 7269 34658 7281 34692
rect 7281 34658 7303 34692
rect 7341 34658 7349 34692
rect 7349 34658 7375 34692
rect 7413 34658 7417 34692
rect 7417 34658 7447 34692
rect 7485 34658 7519 34692
rect 7557 34658 7587 34692
rect 7587 34658 7591 34692
rect 7629 34658 7655 34692
rect 7655 34658 7663 34692
rect 7701 34658 7723 34692
rect 7723 34658 7735 34692
rect 7773 34658 7791 34692
rect 7791 34658 7807 34692
rect 7845 34658 7859 34692
rect 7859 34658 7879 34692
rect 7917 34658 7927 34692
rect 7927 34658 7951 34692
rect 7989 34658 7995 34692
rect 7995 34658 8023 34692
rect 8061 34658 8063 34692
rect 8063 34658 8095 34692
rect 8133 34658 8165 34692
rect 8165 34658 8167 34692
rect 8205 34658 8233 34692
rect 8233 34658 8239 34692
rect 8277 34658 8301 34692
rect 8301 34658 8311 34692
rect 8349 34658 8369 34692
rect 8369 34658 8383 34692
rect 8421 34658 8437 34692
rect 8437 34658 8455 34692
rect 8493 34658 8505 34692
rect 8505 34658 8527 34692
rect 8565 34658 8573 34692
rect 8573 34658 8599 34692
rect 8637 34658 8641 34692
rect 8641 34658 8671 34692
rect 8709 34658 8743 34692
rect 8781 34658 8811 34692
rect 8811 34658 8815 34692
rect 8853 34658 8879 34692
rect 8879 34658 8887 34692
rect 8925 34658 8947 34692
rect 8947 34658 8959 34692
rect 8997 34658 9015 34692
rect 9015 34658 9031 34692
rect 9069 34658 9083 34692
rect 9083 34658 9103 34692
rect 9141 34658 9151 34692
rect 9151 34658 9175 34692
rect 9213 34658 9219 34692
rect 9219 34658 9247 34692
rect 9285 34658 9287 34692
rect 9287 34658 9319 34692
rect 9357 34658 9389 34692
rect 9389 34658 9391 34692
rect 9429 34658 9457 34692
rect 9457 34658 9463 34692
rect 9501 34658 9525 34692
rect 9525 34658 9535 34692
rect 9573 34658 9593 34692
rect 9593 34658 9607 34692
rect 9645 34658 9661 34692
rect 9661 34658 9679 34692
rect 9717 34658 9729 34692
rect 9729 34658 9751 34692
rect 9789 34658 9797 34692
rect 9797 34658 9823 34692
rect 9861 34658 9865 34692
rect 9865 34658 9895 34692
rect 9933 34658 9967 34692
rect 10005 34658 10035 34692
rect 10035 34658 10039 34692
rect 10077 34658 10103 34692
rect 10103 34658 10111 34692
rect 10149 34658 10171 34692
rect 10171 34658 10183 34692
rect 10221 34658 10239 34692
rect 10239 34658 10255 34692
rect 10293 34658 10307 34692
rect 10307 34658 10327 34692
rect 10365 34658 10375 34692
rect 10375 34658 10399 34692
rect 10437 34658 10443 34692
rect 10443 34658 10471 34692
rect 10509 34658 10511 34692
rect 10511 34658 10543 34692
rect 10581 34658 10613 34692
rect 10613 34658 10615 34692
rect 10653 34658 10681 34692
rect 10681 34658 10687 34692
rect 10725 34658 10749 34692
rect 10749 34658 10759 34692
rect 10797 34658 10817 34692
rect 10817 34658 10831 34692
rect 10869 34658 10885 34692
rect 10885 34658 10903 34692
rect 10941 34658 10953 34692
rect 10953 34658 10975 34692
rect 11013 34658 11021 34692
rect 11021 34658 11047 34692
rect 11085 34658 11089 34692
rect 11089 34658 11119 34692
rect 11157 34658 11191 34692
rect 11229 34658 11259 34692
rect 11259 34658 11263 34692
rect 11301 34658 11327 34692
rect 11327 34658 11335 34692
rect 11373 34658 11395 34692
rect 11395 34658 11407 34692
rect 11445 34658 11463 34692
rect 11463 34658 11479 34692
rect 11517 34658 11531 34692
rect 11531 34658 11551 34692
rect 11589 34658 11599 34692
rect 11599 34658 11623 34692
rect 11661 34658 11667 34692
rect 11667 34658 11695 34692
rect 11733 34658 11735 34692
rect 11735 34658 11767 34692
rect 11805 34658 11837 34692
rect 11837 34658 11839 34692
rect 11877 34658 11905 34692
rect 11905 34658 11911 34692
rect 11949 34658 11973 34692
rect 11973 34658 11983 34692
rect 12021 34658 12041 34692
rect 12041 34658 12055 34692
rect 12093 34658 12109 34692
rect 12109 34658 12127 34692
rect 12165 34658 12177 34692
rect 12177 34658 12199 34692
rect 12237 34658 12245 34692
rect 12245 34658 12271 34692
rect 12309 34658 12313 34692
rect 12313 34658 12343 34692
rect 12381 34658 12415 34692
rect 12453 34658 12483 34692
rect 12483 34658 12487 34692
rect 12525 34658 12551 34692
rect 12551 34658 12559 34692
rect 12597 34658 12619 34692
rect 12619 34658 12631 34692
rect 12669 34658 12687 34692
rect 12687 34658 12703 34692
rect 12741 34658 12755 34692
rect 12755 34658 12775 34692
rect 12813 34658 12823 34692
rect 12823 34658 12847 34692
rect 12885 34658 12891 34692
rect 12891 34658 12919 34692
rect 12957 34658 12959 34692
rect 12959 34658 12991 34692
rect 13029 34658 13061 34692
rect 13061 34658 13063 34692
rect 13101 34658 13129 34692
rect 13129 34658 13135 34692
rect 13173 34658 13197 34692
rect 13197 34658 13207 34692
rect 13245 34658 13265 34692
rect 13265 34658 13279 34692
rect 13317 34658 13333 34692
rect 13333 34658 13351 34692
rect 13389 34658 13401 34692
rect 13401 34658 13423 34692
rect 13461 34658 13469 34692
rect 13469 34658 13495 34692
rect 13533 34658 13537 34692
rect 13537 34658 13567 34692
rect 13605 34658 13639 34692
rect 13677 34658 13707 34692
rect 13707 34658 13711 34692
rect 1153 34475 1187 34495
rect 1153 34461 1187 34475
rect 1153 34407 1187 34423
rect 1153 34389 1187 34407
rect 1153 34339 1187 34351
rect 1153 34317 1187 34339
rect 1153 34271 1187 34279
rect 1153 34245 1187 34271
rect 1153 34203 1187 34207
rect 1153 34173 1187 34203
rect 1153 34101 1187 34135
rect 1153 34033 1187 34063
rect 1153 34029 1187 34033
rect 1153 33965 1187 33991
rect 1153 33957 1187 33965
rect 1153 33897 1187 33919
rect 1153 33885 1187 33897
rect 1153 33829 1187 33847
rect 1153 33813 1187 33829
rect 1153 33761 1187 33775
rect 1153 33741 1187 33761
rect 1153 33693 1187 33703
rect 1153 33669 1187 33693
rect 1153 33625 1187 33631
rect 1153 33597 1187 33625
rect 1153 33557 1187 33559
rect 1153 33525 1187 33557
rect 1153 33455 1187 33487
rect 1153 33453 1187 33455
rect 1153 33387 1187 33415
rect 1153 33381 1187 33387
rect 1153 33319 1187 33343
rect 1153 33309 1187 33319
rect 1153 33251 1187 33271
rect 1153 33237 1187 33251
rect 1153 33183 1187 33199
rect 1153 33165 1187 33183
rect 1153 33115 1187 33127
rect 1153 33093 1187 33115
rect 1153 33047 1187 33055
rect 1153 33021 1187 33047
rect 1153 32979 1187 32983
rect 1153 32949 1187 32979
rect 1153 32877 1187 32911
rect 1153 32809 1187 32839
rect 1153 32805 1187 32809
rect 1153 32741 1187 32767
rect 1153 32733 1187 32741
rect 1153 32673 1187 32695
rect 1153 32661 1187 32673
rect 1153 32605 1187 32623
rect 1153 32589 1187 32605
rect 1153 32537 1187 32551
rect 1153 32517 1187 32537
rect 1153 32469 1187 32479
rect 1153 32445 1187 32469
rect 1153 32401 1187 32407
rect 1153 32373 1187 32401
rect 1153 32333 1187 32335
rect 1153 32301 1187 32333
rect 1153 32231 1187 32263
rect 1153 32229 1187 32231
rect 1153 32163 1187 32191
rect 1153 32157 1187 32163
rect 1153 32095 1187 32119
rect 1153 32085 1187 32095
rect 1153 32027 1187 32047
rect 1153 32013 1187 32027
rect 1153 31959 1187 31975
rect 1153 31941 1187 31959
rect 1153 31891 1187 31903
rect 1153 31869 1187 31891
rect 1153 31823 1187 31831
rect 1153 31797 1187 31823
rect 1153 31755 1187 31759
rect 1153 31725 1187 31755
rect 1153 31653 1187 31687
rect 1153 31585 1187 31615
rect 1153 31581 1187 31585
rect 1153 31517 1187 31543
rect 1153 31509 1187 31517
rect 1153 31449 1187 31471
rect 1153 31437 1187 31449
rect 1153 31381 1187 31399
rect 1153 31365 1187 31381
rect 1153 31313 1187 31327
rect 1153 31293 1187 31313
rect 1153 31245 1187 31255
rect 1153 31221 1187 31245
rect 1153 31177 1187 31183
rect 1153 31149 1187 31177
rect 1153 31109 1187 31111
rect 1153 31077 1187 31109
rect 1153 31007 1187 31039
rect 1153 31005 1187 31007
rect 1153 30939 1187 30967
rect 1153 30933 1187 30939
rect 1153 30871 1187 30895
rect 1153 30861 1187 30871
rect 1153 30803 1187 30823
rect 1153 30789 1187 30803
rect 1153 30735 1187 30751
rect 1153 30717 1187 30735
rect 1153 30667 1187 30679
rect 1153 30645 1187 30667
rect 1153 30599 1187 30607
rect 1153 30573 1187 30599
rect 1153 30531 1187 30535
rect 1153 30501 1187 30531
rect 1153 30429 1187 30463
rect 1153 30361 1187 30391
rect 1153 30357 1187 30361
rect 1153 30293 1187 30319
rect 1153 30285 1187 30293
rect 1153 30225 1187 30247
rect 1153 30213 1187 30225
rect 1153 30157 1187 30175
rect 1153 30141 1187 30157
rect 1153 30089 1187 30103
rect 1153 30069 1187 30089
rect 1153 30021 1187 30031
rect 1153 29997 1187 30021
rect 1153 29953 1187 29959
rect 1153 29925 1187 29953
rect 1153 29885 1187 29887
rect 1153 29853 1187 29885
rect 1153 29783 1187 29815
rect 1153 29781 1187 29783
rect 1153 29715 1187 29743
rect 1153 29709 1187 29715
rect 1153 29647 1187 29671
rect 1153 29637 1187 29647
rect 1153 29579 1187 29599
rect 1153 29565 1187 29579
rect 1153 29511 1187 29527
rect 1153 29493 1187 29511
rect 1153 29443 1187 29455
rect 1153 29421 1187 29443
rect 1153 29375 1187 29383
rect 1153 29349 1187 29375
rect 1153 29307 1187 29311
rect 1153 29277 1187 29307
rect 1153 29205 1187 29239
rect 1153 29137 1187 29167
rect 1153 29133 1187 29137
rect 1153 29069 1187 29095
rect 1153 29061 1187 29069
rect 1153 29001 1187 29023
rect 1153 28989 1187 29001
rect 1153 28933 1187 28951
rect 1153 28917 1187 28933
rect 13801 34470 13835 34487
rect 13801 34453 13835 34470
rect 13801 34402 13835 34415
rect 13801 34381 13835 34402
rect 13801 34334 13835 34343
rect 13801 34309 13835 34334
rect 13801 34266 13835 34271
rect 13801 34237 13835 34266
rect 13801 34198 13835 34199
rect 13801 34165 13835 34198
rect 13801 34096 13835 34127
rect 13801 34093 13835 34096
rect 13801 34028 13835 34055
rect 13801 34021 13835 34028
rect 13801 33960 13835 33983
rect 13801 33949 13835 33960
rect 13801 33892 13835 33911
rect 13801 33877 13835 33892
rect 13801 33824 13835 33839
rect 13801 33805 13835 33824
rect 13801 33756 13835 33767
rect 13801 33733 13835 33756
rect 13801 33688 13835 33695
rect 13801 33661 13835 33688
rect 13801 33620 13835 33623
rect 13801 33589 13835 33620
rect 13801 33518 13835 33551
rect 13801 33517 13835 33518
rect 13801 33450 13835 33479
rect 13801 33445 13835 33450
rect 13801 33382 13835 33407
rect 13801 33373 13835 33382
rect 13801 33314 13835 33335
rect 13801 33301 13835 33314
rect 13801 33246 13835 33263
rect 13801 33229 13835 33246
rect 13801 33178 13835 33191
rect 13801 33157 13835 33178
rect 13801 33110 13835 33119
rect 13801 33085 13835 33110
rect 13801 33042 13835 33047
rect 13801 33013 13835 33042
rect 13801 32974 13835 32975
rect 13801 32941 13835 32974
rect 13801 32872 13835 32903
rect 13801 32869 13835 32872
rect 13801 32804 13835 32831
rect 13801 32797 13835 32804
rect 13801 32736 13835 32759
rect 13801 32725 13835 32736
rect 13801 32668 13835 32687
rect 13801 32653 13835 32668
rect 13801 32600 13835 32615
rect 13801 32581 13835 32600
rect 13801 32532 13835 32543
rect 13801 32509 13835 32532
rect 13801 32464 13835 32471
rect 13801 32437 13835 32464
rect 13801 32396 13835 32399
rect 13801 32365 13835 32396
rect 13801 32294 13835 32327
rect 13801 32293 13835 32294
rect 13801 32226 13835 32255
rect 13801 32221 13835 32226
rect 13801 32158 13835 32183
rect 13801 32149 13835 32158
rect 13801 32090 13835 32111
rect 13801 32077 13835 32090
rect 13801 32022 13835 32039
rect 13801 32005 13835 32022
rect 13801 31954 13835 31967
rect 13801 31933 13835 31954
rect 13801 31886 13835 31895
rect 13801 31861 13835 31886
rect 13801 31818 13835 31823
rect 13801 31789 13835 31818
rect 13801 31750 13835 31751
rect 13801 31717 13835 31750
rect 13801 31648 13835 31679
rect 13801 31645 13835 31648
rect 13801 31580 13835 31607
rect 13801 31573 13835 31580
rect 13801 31512 13835 31535
rect 13801 31501 13835 31512
rect 13801 31444 13835 31463
rect 13801 31429 13835 31444
rect 13801 31376 13835 31391
rect 13801 31357 13835 31376
rect 13801 31308 13835 31319
rect 13801 31285 13835 31308
rect 13801 31240 13835 31247
rect 13801 31213 13835 31240
rect 13801 31172 13835 31175
rect 13801 31141 13835 31172
rect 13801 31070 13835 31103
rect 13801 31069 13835 31070
rect 13801 31002 13835 31031
rect 13801 30997 13835 31002
rect 13801 30934 13835 30959
rect 13801 30925 13835 30934
rect 13801 30866 13835 30887
rect 13801 30853 13835 30866
rect 13801 30798 13835 30815
rect 13801 30781 13835 30798
rect 13801 30730 13835 30743
rect 13801 30709 13835 30730
rect 13801 30662 13835 30671
rect 13801 30637 13835 30662
rect 13801 30594 13835 30599
rect 13801 30565 13835 30594
rect 13801 30526 13835 30527
rect 13801 30493 13835 30526
rect 13801 30424 13835 30455
rect 13801 30421 13835 30424
rect 13801 30356 13835 30383
rect 13801 30349 13835 30356
rect 13801 30288 13835 30311
rect 13801 30277 13835 30288
rect 13801 30220 13835 30239
rect 13801 30205 13835 30220
rect 13801 30152 13835 30167
rect 13801 30133 13835 30152
rect 13801 30084 13835 30095
rect 13801 30061 13835 30084
rect 13801 30016 13835 30023
rect 13801 29989 13835 30016
rect 13801 29948 13835 29951
rect 13801 29917 13835 29948
rect 13801 29846 13835 29879
rect 13801 29845 13835 29846
rect 13801 29778 13835 29807
rect 13801 29773 13835 29778
rect 13801 29710 13835 29735
rect 13801 29701 13835 29710
rect 13801 29642 13835 29663
rect 13801 29629 13835 29642
rect 13801 29574 13835 29591
rect 13801 29557 13835 29574
rect 13801 29506 13835 29519
rect 13801 29485 13835 29506
rect 13801 29438 13835 29447
rect 13801 29413 13835 29438
rect 13801 29370 13835 29375
rect 13801 29341 13835 29370
rect 13801 29302 13835 29303
rect 13801 29269 13835 29302
rect 13801 29200 13835 29231
rect 13801 29197 13835 29200
rect 13801 29132 13835 29159
rect 13801 29125 13835 29132
rect 13801 29064 13835 29087
rect 13801 29053 13835 29064
rect 13801 28996 13835 29015
rect 13801 28981 13835 28996
rect 1153 28865 1187 28879
rect 1153 28845 1187 28865
rect 1153 28797 1187 28807
rect 1153 28773 1187 28797
rect 1153 28729 1187 28735
rect 1153 28701 1187 28729
rect 1153 28661 1187 28663
rect 1153 28629 1187 28661
rect 1153 28559 1187 28591
rect 1153 28557 1187 28559
rect 1153 28491 1187 28519
rect 1153 28485 1187 28491
rect 1153 28423 1187 28447
rect 1153 28413 1187 28423
rect 1153 28355 1187 28375
rect 1153 28341 1187 28355
rect 1153 28287 1187 28303
rect 1153 28269 1187 28287
rect 1153 28219 1187 28231
rect 1153 28197 1187 28219
rect 1153 28151 1187 28159
rect 1153 28125 1187 28151
rect 1153 28083 1187 28087
rect 1153 28053 1187 28083
rect 1153 27981 1187 28015
rect 1153 27913 1187 27943
rect 1153 27909 1187 27913
rect 1153 27845 1187 27871
rect 1153 27837 1187 27845
rect 1153 27777 1187 27799
rect 1153 27765 1187 27777
rect 1153 27709 1187 27727
rect 1153 27693 1187 27709
rect 1153 27641 1187 27655
rect 1153 27621 1187 27641
rect 1153 27573 1187 27583
rect 1153 27549 1187 27573
rect 1153 27505 1187 27511
rect 1153 27477 1187 27505
rect 1153 27437 1187 27439
rect 1153 27405 1187 27437
rect 1153 27335 1187 27367
rect 1153 27333 1187 27335
rect 1153 27267 1187 27295
rect 1153 27261 1187 27267
rect 1153 27199 1187 27223
rect 1153 27189 1187 27199
rect 1153 27131 1187 27151
rect 1153 27117 1187 27131
rect 1153 27063 1187 27079
rect 1153 27045 1187 27063
rect 1974 28566 2111 28888
rect 2111 28566 12889 28888
rect 12889 28566 13024 28888
rect 1718 28435 1968 28502
rect 1718 27517 1968 28435
rect 13023 28435 13273 28495
rect 2443 28243 2477 28277
rect 2515 28273 2549 28277
rect 2515 28243 2519 28273
rect 2519 28243 2549 28273
rect 2587 28243 2621 28277
rect 2659 28273 2693 28277
rect 2731 28273 2765 28277
rect 2803 28273 2837 28277
rect 2875 28273 2909 28277
rect 2947 28273 2981 28277
rect 3019 28273 3053 28277
rect 3091 28273 3125 28277
rect 3163 28273 3197 28277
rect 3235 28273 3269 28277
rect 3307 28273 3341 28277
rect 3379 28273 3413 28277
rect 3451 28273 3485 28277
rect 3523 28273 3557 28277
rect 3595 28273 3629 28277
rect 3667 28273 3701 28277
rect 3739 28273 3773 28277
rect 2659 28243 2689 28273
rect 2689 28243 2693 28273
rect 2731 28243 2757 28273
rect 2757 28243 2765 28273
rect 2803 28243 2825 28273
rect 2825 28243 2837 28273
rect 2875 28243 2893 28273
rect 2893 28243 2909 28273
rect 2947 28243 2961 28273
rect 2961 28243 2981 28273
rect 3019 28243 3029 28273
rect 3029 28243 3053 28273
rect 3091 28243 3097 28273
rect 3097 28243 3125 28273
rect 3163 28243 3165 28273
rect 3165 28243 3197 28273
rect 3235 28243 3267 28273
rect 3267 28243 3269 28273
rect 3307 28243 3335 28273
rect 3335 28243 3341 28273
rect 3379 28243 3403 28273
rect 3403 28243 3413 28273
rect 3451 28243 3471 28273
rect 3471 28243 3485 28273
rect 3523 28243 3539 28273
rect 3539 28243 3557 28273
rect 3595 28243 3607 28273
rect 3607 28243 3629 28273
rect 3667 28243 3675 28273
rect 3675 28243 3701 28273
rect 3739 28243 3743 28273
rect 3743 28243 3773 28273
rect 3811 28243 3845 28277
rect 3883 28273 3917 28277
rect 3955 28273 3989 28277
rect 4027 28273 4061 28277
rect 4099 28273 4133 28277
rect 4171 28273 4205 28277
rect 4243 28273 4277 28277
rect 4315 28273 4349 28277
rect 4387 28273 4421 28277
rect 4459 28273 4493 28277
rect 4531 28273 4565 28277
rect 4603 28273 4637 28277
rect 4675 28273 4709 28277
rect 4747 28273 4781 28277
rect 4819 28273 4853 28277
rect 4891 28273 4925 28277
rect 4963 28273 4997 28277
rect 3883 28243 3913 28273
rect 3913 28243 3917 28273
rect 3955 28243 3981 28273
rect 3981 28243 3989 28273
rect 4027 28243 4049 28273
rect 4049 28243 4061 28273
rect 4099 28243 4117 28273
rect 4117 28243 4133 28273
rect 4171 28243 4185 28273
rect 4185 28243 4205 28273
rect 4243 28243 4253 28273
rect 4253 28243 4277 28273
rect 4315 28243 4321 28273
rect 4321 28243 4349 28273
rect 4387 28243 4389 28273
rect 4389 28243 4421 28273
rect 4459 28243 4491 28273
rect 4491 28243 4493 28273
rect 4531 28243 4559 28273
rect 4559 28243 4565 28273
rect 4603 28243 4627 28273
rect 4627 28243 4637 28273
rect 4675 28243 4695 28273
rect 4695 28243 4709 28273
rect 4747 28243 4763 28273
rect 4763 28243 4781 28273
rect 4819 28243 4831 28273
rect 4831 28243 4853 28273
rect 4891 28243 4899 28273
rect 4899 28243 4925 28273
rect 4963 28243 4967 28273
rect 4967 28243 4997 28273
rect 5035 28243 5069 28277
rect 5107 28273 5141 28277
rect 5179 28273 5213 28277
rect 5251 28273 5285 28277
rect 5323 28273 5357 28277
rect 5395 28273 5429 28277
rect 5467 28273 5501 28277
rect 5539 28273 5573 28277
rect 5611 28273 5645 28277
rect 5683 28273 5717 28277
rect 5755 28273 5789 28277
rect 5827 28273 5861 28277
rect 5899 28273 5933 28277
rect 5971 28273 6005 28277
rect 6043 28273 6077 28277
rect 6115 28273 6149 28277
rect 6187 28273 6221 28277
rect 5107 28243 5137 28273
rect 5137 28243 5141 28273
rect 5179 28243 5205 28273
rect 5205 28243 5213 28273
rect 5251 28243 5273 28273
rect 5273 28243 5285 28273
rect 5323 28243 5341 28273
rect 5341 28243 5357 28273
rect 5395 28243 5409 28273
rect 5409 28243 5429 28273
rect 5467 28243 5477 28273
rect 5477 28243 5501 28273
rect 5539 28243 5545 28273
rect 5545 28243 5573 28273
rect 5611 28243 5613 28273
rect 5613 28243 5645 28273
rect 5683 28243 5715 28273
rect 5715 28243 5717 28273
rect 5755 28243 5783 28273
rect 5783 28243 5789 28273
rect 5827 28243 5851 28273
rect 5851 28243 5861 28273
rect 5899 28243 5919 28273
rect 5919 28243 5933 28273
rect 5971 28243 5987 28273
rect 5987 28243 6005 28273
rect 6043 28243 6055 28273
rect 6055 28243 6077 28273
rect 6115 28243 6123 28273
rect 6123 28243 6149 28273
rect 6187 28243 6191 28273
rect 6191 28243 6221 28273
rect 6259 28243 6293 28277
rect 6331 28273 6365 28277
rect 6403 28273 6437 28277
rect 6475 28273 6509 28277
rect 6547 28273 6581 28277
rect 6619 28273 6653 28277
rect 6691 28273 6725 28277
rect 6763 28273 6797 28277
rect 6835 28273 6869 28277
rect 6907 28273 6941 28277
rect 6979 28273 7013 28277
rect 7051 28273 7085 28277
rect 7123 28273 7157 28277
rect 7195 28273 7229 28277
rect 7267 28273 7301 28277
rect 7339 28273 7373 28277
rect 7411 28273 7445 28277
rect 6331 28243 6361 28273
rect 6361 28243 6365 28273
rect 6403 28243 6429 28273
rect 6429 28243 6437 28273
rect 6475 28243 6497 28273
rect 6497 28243 6509 28273
rect 6547 28243 6565 28273
rect 6565 28243 6581 28273
rect 6619 28243 6633 28273
rect 6633 28243 6653 28273
rect 6691 28243 6701 28273
rect 6701 28243 6725 28273
rect 6763 28243 6769 28273
rect 6769 28243 6797 28273
rect 6835 28243 6837 28273
rect 6837 28243 6869 28273
rect 6907 28243 6939 28273
rect 6939 28243 6941 28273
rect 6979 28243 7007 28273
rect 7007 28243 7013 28273
rect 7051 28243 7075 28273
rect 7075 28243 7085 28273
rect 7123 28243 7143 28273
rect 7143 28243 7157 28273
rect 7195 28243 7211 28273
rect 7211 28243 7229 28273
rect 7267 28243 7279 28273
rect 7279 28243 7301 28273
rect 7339 28243 7347 28273
rect 7347 28243 7373 28273
rect 7411 28243 7415 28273
rect 7415 28243 7445 28273
rect 7483 28243 7517 28277
rect 7555 28273 7589 28277
rect 7627 28273 7661 28277
rect 7699 28273 7733 28277
rect 7771 28273 7805 28277
rect 7843 28273 7877 28277
rect 7915 28273 7949 28277
rect 7987 28273 8021 28277
rect 8059 28273 8093 28277
rect 8131 28273 8165 28277
rect 8203 28273 8237 28277
rect 8275 28273 8309 28277
rect 8347 28273 8381 28277
rect 8419 28273 8453 28277
rect 8491 28273 8525 28277
rect 8563 28273 8597 28277
rect 8635 28273 8669 28277
rect 7555 28243 7585 28273
rect 7585 28243 7589 28273
rect 7627 28243 7653 28273
rect 7653 28243 7661 28273
rect 7699 28243 7721 28273
rect 7721 28243 7733 28273
rect 7771 28243 7789 28273
rect 7789 28243 7805 28273
rect 7843 28243 7857 28273
rect 7857 28243 7877 28273
rect 7915 28243 7925 28273
rect 7925 28243 7949 28273
rect 7987 28243 7993 28273
rect 7993 28243 8021 28273
rect 8059 28243 8061 28273
rect 8061 28243 8093 28273
rect 8131 28243 8163 28273
rect 8163 28243 8165 28273
rect 8203 28243 8231 28273
rect 8231 28243 8237 28273
rect 8275 28243 8299 28273
rect 8299 28243 8309 28273
rect 8347 28243 8367 28273
rect 8367 28243 8381 28273
rect 8419 28243 8435 28273
rect 8435 28243 8453 28273
rect 8491 28243 8503 28273
rect 8503 28243 8525 28273
rect 8563 28243 8571 28273
rect 8571 28243 8597 28273
rect 8635 28243 8639 28273
rect 8639 28243 8669 28273
rect 8707 28243 8741 28277
rect 8779 28273 8813 28277
rect 8851 28273 8885 28277
rect 8923 28273 8957 28277
rect 8995 28273 9029 28277
rect 9067 28273 9101 28277
rect 9139 28273 9173 28277
rect 9211 28273 9245 28277
rect 9283 28273 9317 28277
rect 9355 28273 9389 28277
rect 9427 28273 9461 28277
rect 9499 28273 9533 28277
rect 9571 28273 9605 28277
rect 9643 28273 9677 28277
rect 9715 28273 9749 28277
rect 9787 28273 9821 28277
rect 9859 28273 9893 28277
rect 8779 28243 8809 28273
rect 8809 28243 8813 28273
rect 8851 28243 8877 28273
rect 8877 28243 8885 28273
rect 8923 28243 8945 28273
rect 8945 28243 8957 28273
rect 8995 28243 9013 28273
rect 9013 28243 9029 28273
rect 9067 28243 9081 28273
rect 9081 28243 9101 28273
rect 9139 28243 9149 28273
rect 9149 28243 9173 28273
rect 9211 28243 9217 28273
rect 9217 28243 9245 28273
rect 9283 28243 9285 28273
rect 9285 28243 9317 28273
rect 9355 28243 9387 28273
rect 9387 28243 9389 28273
rect 9427 28243 9455 28273
rect 9455 28243 9461 28273
rect 9499 28243 9523 28273
rect 9523 28243 9533 28273
rect 9571 28243 9591 28273
rect 9591 28243 9605 28273
rect 9643 28243 9659 28273
rect 9659 28243 9677 28273
rect 9715 28243 9727 28273
rect 9727 28243 9749 28273
rect 9787 28243 9795 28273
rect 9795 28243 9821 28273
rect 9859 28243 9863 28273
rect 9863 28243 9893 28273
rect 9931 28243 9965 28277
rect 10003 28273 10037 28277
rect 10075 28273 10109 28277
rect 10147 28273 10181 28277
rect 10219 28273 10253 28277
rect 10291 28273 10325 28277
rect 10363 28273 10397 28277
rect 10435 28273 10469 28277
rect 10507 28273 10541 28277
rect 10579 28273 10613 28277
rect 10651 28273 10685 28277
rect 10723 28273 10757 28277
rect 10795 28273 10829 28277
rect 10867 28273 10901 28277
rect 10939 28273 10973 28277
rect 11011 28273 11045 28277
rect 11083 28273 11117 28277
rect 10003 28243 10033 28273
rect 10033 28243 10037 28273
rect 10075 28243 10101 28273
rect 10101 28243 10109 28273
rect 10147 28243 10169 28273
rect 10169 28243 10181 28273
rect 10219 28243 10237 28273
rect 10237 28243 10253 28273
rect 10291 28243 10305 28273
rect 10305 28243 10325 28273
rect 10363 28243 10373 28273
rect 10373 28243 10397 28273
rect 10435 28243 10441 28273
rect 10441 28243 10469 28273
rect 10507 28243 10509 28273
rect 10509 28243 10541 28273
rect 10579 28243 10611 28273
rect 10611 28243 10613 28273
rect 10651 28243 10679 28273
rect 10679 28243 10685 28273
rect 10723 28243 10747 28273
rect 10747 28243 10757 28273
rect 10795 28243 10815 28273
rect 10815 28243 10829 28273
rect 10867 28243 10883 28273
rect 10883 28243 10901 28273
rect 10939 28243 10951 28273
rect 10951 28243 10973 28273
rect 11011 28243 11019 28273
rect 11019 28243 11045 28273
rect 11083 28243 11087 28273
rect 11087 28243 11117 28273
rect 11155 28243 11189 28277
rect 11227 28273 11261 28277
rect 11299 28273 11333 28277
rect 11371 28273 11405 28277
rect 11443 28273 11477 28277
rect 11515 28273 11549 28277
rect 11587 28273 11621 28277
rect 11659 28273 11693 28277
rect 11731 28273 11765 28277
rect 11803 28273 11837 28277
rect 11875 28273 11909 28277
rect 11947 28273 11981 28277
rect 12019 28273 12053 28277
rect 12091 28273 12125 28277
rect 12163 28273 12197 28277
rect 12235 28273 12269 28277
rect 12307 28273 12341 28277
rect 11227 28243 11257 28273
rect 11257 28243 11261 28273
rect 11299 28243 11325 28273
rect 11325 28243 11333 28273
rect 11371 28243 11393 28273
rect 11393 28243 11405 28273
rect 11443 28243 11461 28273
rect 11461 28243 11477 28273
rect 11515 28243 11529 28273
rect 11529 28243 11549 28273
rect 11587 28243 11597 28273
rect 11597 28243 11621 28273
rect 11659 28243 11665 28273
rect 11665 28243 11693 28273
rect 11731 28243 11733 28273
rect 11733 28243 11765 28273
rect 11803 28243 11835 28273
rect 11835 28243 11837 28273
rect 11875 28243 11903 28273
rect 11903 28243 11909 28273
rect 11947 28243 11971 28273
rect 11971 28243 11981 28273
rect 12019 28243 12039 28273
rect 12039 28243 12053 28273
rect 12091 28243 12107 28273
rect 12107 28243 12125 28273
rect 12163 28243 12175 28273
rect 12175 28243 12197 28273
rect 12235 28243 12243 28273
rect 12243 28243 12269 28273
rect 12307 28243 12311 28273
rect 12311 28243 12341 28273
rect 12379 28243 12413 28277
rect 12451 28273 12485 28277
rect 12451 28243 12481 28273
rect 12481 28243 12485 28273
rect 12523 28243 12557 28277
rect 2479 28169 2485 28203
rect 2485 28169 2513 28203
rect 2551 28169 2553 28203
rect 2553 28169 2585 28203
rect 2623 28169 2655 28203
rect 2655 28169 2657 28203
rect 2695 28169 2723 28203
rect 2723 28169 2729 28203
rect 2767 28169 2791 28203
rect 2791 28169 2801 28203
rect 2839 28169 2859 28203
rect 2859 28169 2873 28203
rect 2911 28169 2927 28203
rect 2927 28169 2945 28203
rect 2983 28169 2995 28203
rect 2995 28169 3017 28203
rect 3055 28169 3063 28203
rect 3063 28169 3089 28203
rect 3127 28169 3131 28203
rect 3131 28169 3161 28203
rect 3199 28169 3233 28203
rect 3271 28169 3301 28203
rect 3301 28169 3305 28203
rect 3343 28169 3369 28203
rect 3369 28169 3377 28203
rect 3415 28169 3437 28203
rect 3437 28169 3449 28203
rect 3487 28169 3505 28203
rect 3505 28169 3521 28203
rect 3559 28169 3573 28203
rect 3573 28169 3593 28203
rect 3631 28169 3641 28203
rect 3641 28169 3665 28203
rect 3703 28169 3709 28203
rect 3709 28169 3737 28203
rect 3775 28169 3777 28203
rect 3777 28169 3809 28203
rect 3847 28169 3879 28203
rect 3879 28169 3881 28203
rect 3919 28169 3947 28203
rect 3947 28169 3953 28203
rect 3991 28169 4015 28203
rect 4015 28169 4025 28203
rect 4063 28169 4083 28203
rect 4083 28169 4097 28203
rect 4135 28169 4151 28203
rect 4151 28169 4169 28203
rect 4207 28169 4219 28203
rect 4219 28169 4241 28203
rect 4279 28169 4287 28203
rect 4287 28169 4313 28203
rect 4351 28169 4355 28203
rect 4355 28169 4385 28203
rect 4423 28169 4457 28203
rect 4495 28169 4525 28203
rect 4525 28169 4529 28203
rect 4567 28169 4593 28203
rect 4593 28169 4601 28203
rect 4639 28169 4661 28203
rect 4661 28169 4673 28203
rect 4711 28169 4729 28203
rect 4729 28169 4745 28203
rect 4783 28169 4797 28203
rect 4797 28169 4817 28203
rect 4855 28169 4865 28203
rect 4865 28169 4889 28203
rect 4927 28169 4933 28203
rect 4933 28169 4961 28203
rect 4999 28169 5001 28203
rect 5001 28169 5033 28203
rect 5071 28169 5103 28203
rect 5103 28169 5105 28203
rect 5143 28169 5171 28203
rect 5171 28169 5177 28203
rect 5215 28169 5239 28203
rect 5239 28169 5249 28203
rect 5287 28169 5307 28203
rect 5307 28169 5321 28203
rect 5359 28169 5375 28203
rect 5375 28169 5393 28203
rect 5431 28169 5443 28203
rect 5443 28169 5465 28203
rect 5503 28169 5511 28203
rect 5511 28169 5537 28203
rect 5575 28169 5579 28203
rect 5579 28169 5609 28203
rect 5647 28169 5681 28203
rect 5719 28169 5749 28203
rect 5749 28169 5753 28203
rect 5791 28169 5817 28203
rect 5817 28169 5825 28203
rect 5863 28169 5885 28203
rect 5885 28169 5897 28203
rect 5935 28169 5953 28203
rect 5953 28169 5969 28203
rect 6007 28169 6021 28203
rect 6021 28169 6041 28203
rect 6079 28169 6089 28203
rect 6089 28169 6113 28203
rect 6151 28169 6157 28203
rect 6157 28169 6185 28203
rect 6223 28169 6225 28203
rect 6225 28169 6257 28203
rect 6295 28169 6327 28203
rect 6327 28169 6329 28203
rect 6367 28169 6395 28203
rect 6395 28169 6401 28203
rect 6439 28169 6463 28203
rect 6463 28169 6473 28203
rect 6511 28169 6531 28203
rect 6531 28169 6545 28203
rect 6583 28169 6599 28203
rect 6599 28169 6617 28203
rect 6655 28169 6667 28203
rect 6667 28169 6689 28203
rect 6727 28169 6735 28203
rect 6735 28169 6761 28203
rect 6799 28169 6803 28203
rect 6803 28169 6833 28203
rect 6871 28169 6905 28203
rect 6943 28169 6973 28203
rect 6973 28169 6977 28203
rect 7015 28169 7041 28203
rect 7041 28169 7049 28203
rect 7087 28169 7109 28203
rect 7109 28169 7121 28203
rect 7159 28169 7177 28203
rect 7177 28169 7193 28203
rect 7231 28169 7245 28203
rect 7245 28169 7265 28203
rect 7303 28169 7313 28203
rect 7313 28169 7337 28203
rect 7375 28169 7381 28203
rect 7381 28169 7409 28203
rect 7447 28169 7449 28203
rect 7449 28169 7481 28203
rect 7519 28169 7551 28203
rect 7551 28169 7553 28203
rect 7591 28169 7619 28203
rect 7619 28169 7625 28203
rect 7663 28169 7687 28203
rect 7687 28169 7697 28203
rect 7735 28169 7755 28203
rect 7755 28169 7769 28203
rect 7807 28169 7823 28203
rect 7823 28169 7841 28203
rect 7879 28169 7891 28203
rect 7891 28169 7913 28203
rect 7951 28169 7959 28203
rect 7959 28169 7985 28203
rect 8023 28169 8027 28203
rect 8027 28169 8057 28203
rect 8095 28169 8129 28203
rect 8167 28169 8197 28203
rect 8197 28169 8201 28203
rect 8239 28169 8265 28203
rect 8265 28169 8273 28203
rect 8311 28169 8333 28203
rect 8333 28169 8345 28203
rect 8383 28169 8401 28203
rect 8401 28169 8417 28203
rect 8455 28169 8469 28203
rect 8469 28169 8489 28203
rect 8527 28169 8537 28203
rect 8537 28169 8561 28203
rect 8599 28169 8605 28203
rect 8605 28169 8633 28203
rect 8671 28169 8673 28203
rect 8673 28169 8705 28203
rect 8743 28169 8775 28203
rect 8775 28169 8777 28203
rect 8815 28169 8843 28203
rect 8843 28169 8849 28203
rect 8887 28169 8911 28203
rect 8911 28169 8921 28203
rect 8959 28169 8979 28203
rect 8979 28169 8993 28203
rect 9031 28169 9047 28203
rect 9047 28169 9065 28203
rect 9103 28169 9115 28203
rect 9115 28169 9137 28203
rect 9175 28169 9183 28203
rect 9183 28169 9209 28203
rect 9247 28169 9251 28203
rect 9251 28169 9281 28203
rect 9319 28169 9353 28203
rect 9391 28169 9421 28203
rect 9421 28169 9425 28203
rect 9463 28169 9489 28203
rect 9489 28169 9497 28203
rect 9535 28169 9557 28203
rect 9557 28169 9569 28203
rect 9607 28169 9625 28203
rect 9625 28169 9641 28203
rect 9679 28169 9693 28203
rect 9693 28169 9713 28203
rect 9751 28169 9761 28203
rect 9761 28169 9785 28203
rect 9823 28169 9829 28203
rect 9829 28169 9857 28203
rect 9895 28169 9897 28203
rect 9897 28169 9929 28203
rect 9967 28169 9999 28203
rect 9999 28169 10001 28203
rect 10039 28169 10067 28203
rect 10067 28169 10073 28203
rect 10111 28169 10135 28203
rect 10135 28169 10145 28203
rect 10183 28169 10203 28203
rect 10203 28169 10217 28203
rect 10255 28169 10271 28203
rect 10271 28169 10289 28203
rect 10327 28169 10339 28203
rect 10339 28169 10361 28203
rect 10399 28169 10407 28203
rect 10407 28169 10433 28203
rect 10471 28169 10475 28203
rect 10475 28169 10505 28203
rect 10543 28169 10577 28203
rect 10615 28169 10645 28203
rect 10645 28169 10649 28203
rect 10687 28169 10713 28203
rect 10713 28169 10721 28203
rect 10759 28169 10781 28203
rect 10781 28169 10793 28203
rect 10831 28169 10849 28203
rect 10849 28169 10865 28203
rect 10903 28169 10917 28203
rect 10917 28169 10937 28203
rect 10975 28169 10985 28203
rect 10985 28169 11009 28203
rect 11047 28169 11053 28203
rect 11053 28169 11081 28203
rect 11119 28169 11121 28203
rect 11121 28169 11153 28203
rect 11191 28169 11223 28203
rect 11223 28169 11225 28203
rect 11263 28169 11291 28203
rect 11291 28169 11297 28203
rect 11335 28169 11359 28203
rect 11359 28169 11369 28203
rect 11407 28169 11427 28203
rect 11427 28169 11441 28203
rect 11479 28169 11495 28203
rect 11495 28169 11513 28203
rect 11551 28169 11563 28203
rect 11563 28169 11585 28203
rect 11623 28169 11631 28203
rect 11631 28169 11657 28203
rect 11695 28169 11699 28203
rect 11699 28169 11729 28203
rect 11767 28169 11801 28203
rect 11839 28169 11869 28203
rect 11869 28169 11873 28203
rect 11911 28169 11937 28203
rect 11937 28169 11945 28203
rect 11983 28169 12005 28203
rect 12005 28169 12017 28203
rect 12055 28169 12073 28203
rect 12073 28169 12089 28203
rect 12127 28169 12141 28203
rect 12141 28169 12161 28203
rect 12199 28169 12209 28203
rect 12209 28169 12233 28203
rect 12271 28169 12277 28203
rect 12277 28169 12305 28203
rect 12343 28169 12345 28203
rect 12345 28169 12377 28203
rect 12415 28169 12447 28203
rect 12447 28169 12449 28203
rect 12487 28169 12515 28203
rect 12515 28169 12521 28203
rect 2376 28098 2410 28104
rect 2376 28070 2410 28098
rect 12590 28098 12624 28104
rect 12590 28070 12624 28098
rect 2376 28030 2410 28032
rect 2376 27998 2410 28030
rect 2376 27928 2410 27960
rect 2376 27926 2410 27928
rect 2515 27926 2519 28032
rect 2519 27926 12481 28032
rect 12481 27926 12485 28032
rect 12590 28030 12624 28032
rect 12590 27998 12624 28030
rect 12590 27928 12624 27960
rect 12590 27926 12624 27928
rect 2376 27860 2410 27888
rect 2376 27854 2410 27860
rect 12590 27860 12624 27888
rect 12590 27854 12624 27860
rect 2443 27683 2477 27717
rect 2479 27687 2485 27789
rect 2485 27687 12515 27789
rect 12515 27687 12521 27789
rect 2479 27683 12521 27687
rect 12523 27683 12557 27717
rect 1718 27460 1968 27517
rect 13023 27517 13273 28435
rect 13023 27453 13273 27517
rect 1977 27097 2111 27347
rect 2111 27097 12889 27347
rect 12889 27097 13027 27347
rect 13801 28928 13835 28943
rect 13801 28909 13835 28928
rect 13801 28860 13835 28871
rect 13801 28837 13835 28860
rect 13801 28792 13835 28799
rect 13801 28765 13835 28792
rect 1153 26995 1187 27007
rect 1153 26973 1187 26995
rect 1153 26927 1187 26935
rect 1153 26901 1187 26927
rect 1153 26859 1187 26863
rect 1153 26829 1187 26859
rect 1153 26757 1187 26791
rect 1153 26689 1187 26719
rect 1153 26685 1187 26689
rect 1153 26621 1187 26647
rect 1153 26613 1187 26621
rect 1153 26553 1187 26575
rect 1153 26541 1187 26553
rect 1153 26485 1187 26503
rect 1153 26469 1187 26485
rect 1153 26417 1187 26431
rect 1153 26397 1187 26417
rect 1153 26349 1187 26359
rect 1153 26325 1187 26349
rect 1153 26281 1187 26287
rect 1153 26253 1187 26281
rect 1153 26213 1187 26215
rect 1153 26181 1187 26213
rect 1153 26111 1187 26143
rect 1153 26109 1187 26111
rect 1153 26043 1187 26071
rect 1153 26037 1187 26043
rect 1153 25975 1187 25999
rect 1153 25965 1187 25975
rect 1153 25907 1187 25927
rect 1153 25893 1187 25907
rect 1153 25839 1187 25855
rect 1153 25821 1187 25839
rect 1153 25771 1187 25783
rect 1153 25749 1187 25771
rect 1153 25703 1187 25711
rect 1153 25677 1187 25703
rect 1153 25635 1187 25639
rect 1153 25605 1187 25635
rect 1153 25533 1187 25567
rect 1153 25465 1187 25495
rect 1153 25461 1187 25465
rect 1153 25397 1187 25423
rect 1153 25389 1187 25397
rect 1153 25329 1187 25351
rect 1153 25317 1187 25329
rect 1153 25261 1187 25279
rect 1153 25245 1187 25261
rect 1153 25193 1187 25207
rect 1153 25173 1187 25193
rect 1153 25125 1187 25135
rect 1153 25101 1187 25125
rect 1153 25057 1187 25063
rect 1153 25029 1187 25057
rect 1153 24989 1187 24991
rect 1153 24957 1187 24989
rect 1153 24887 1187 24919
rect 1153 24885 1187 24887
rect 1153 24819 1187 24847
rect 1153 24813 1187 24819
rect 2251 26575 12725 26585
rect 2251 26201 2269 26575
rect 2269 26201 12707 26575
rect 12707 26201 12725 26575
rect 2251 26191 12725 26201
rect 1748 26067 2142 26087
rect 1748 25353 1758 26067
rect 1758 25353 2132 26067
rect 2132 25353 2142 26067
rect 1748 25333 2142 25353
rect 2503 25875 2507 25909
rect 2507 25875 2537 25909
rect 2575 25875 2609 25909
rect 2647 25875 2677 25909
rect 2677 25875 2681 25909
rect 2719 25875 2745 25909
rect 2745 25875 2753 25909
rect 2791 25875 2813 25909
rect 2813 25875 2825 25909
rect 2863 25875 2881 25909
rect 2881 25875 2897 25909
rect 2935 25875 2949 25909
rect 2949 25875 2969 25909
rect 3007 25875 3017 25909
rect 3017 25875 3041 25909
rect 3079 25875 3085 25909
rect 3085 25875 3113 25909
rect 3151 25875 3153 25909
rect 3153 25875 3185 25909
rect 3223 25875 3255 25909
rect 3255 25875 3257 25909
rect 3295 25875 3323 25909
rect 3323 25875 3329 25909
rect 3367 25875 3391 25909
rect 3391 25875 3401 25909
rect 3439 25875 3459 25909
rect 3459 25875 3473 25909
rect 3511 25875 3527 25909
rect 3527 25875 3545 25909
rect 3583 25875 3595 25909
rect 3595 25875 3617 25909
rect 3655 25875 3663 25909
rect 3663 25875 3689 25909
rect 3727 25875 3731 25909
rect 3731 25875 3761 25909
rect 3799 25875 3833 25909
rect 3871 25875 3901 25909
rect 3901 25875 3905 25909
rect 3943 25875 3969 25909
rect 3969 25875 3977 25909
rect 4015 25875 4037 25909
rect 4037 25875 4049 25909
rect 4087 25875 4105 25909
rect 4105 25875 4121 25909
rect 4159 25875 4173 25909
rect 4173 25875 4193 25909
rect 4231 25875 4241 25909
rect 4241 25875 4265 25909
rect 4303 25875 4309 25909
rect 4309 25875 4337 25909
rect 4375 25875 4377 25909
rect 4377 25875 4409 25909
rect 4447 25875 4479 25909
rect 4479 25875 4481 25909
rect 4519 25875 4547 25909
rect 4547 25875 4553 25909
rect 4591 25875 4615 25909
rect 4615 25875 4625 25909
rect 4663 25875 4683 25909
rect 4683 25875 4697 25909
rect 4735 25875 4751 25909
rect 4751 25875 4769 25909
rect 4807 25875 4819 25909
rect 4819 25875 4841 25909
rect 4879 25875 4887 25909
rect 4887 25875 4913 25909
rect 4951 25875 4955 25909
rect 4955 25875 4985 25909
rect 5023 25875 5057 25909
rect 5095 25875 5125 25909
rect 5125 25875 5129 25909
rect 5167 25875 5193 25909
rect 5193 25875 5201 25909
rect 5239 25875 5261 25909
rect 5261 25875 5273 25909
rect 5311 25875 5329 25909
rect 5329 25875 5345 25909
rect 5383 25875 5397 25909
rect 5397 25875 5417 25909
rect 5455 25875 5465 25909
rect 5465 25875 5489 25909
rect 5527 25875 5533 25909
rect 5533 25875 5561 25909
rect 5599 25875 5601 25909
rect 5601 25875 5633 25909
rect 5671 25875 5703 25909
rect 5703 25875 5705 25909
rect 5743 25875 5771 25909
rect 5771 25875 5777 25909
rect 5815 25875 5839 25909
rect 5839 25875 5849 25909
rect 5887 25875 5907 25909
rect 5907 25875 5921 25909
rect 5959 25875 5975 25909
rect 5975 25875 5993 25909
rect 6031 25875 6043 25909
rect 6043 25875 6065 25909
rect 6103 25875 6111 25909
rect 6111 25875 6137 25909
rect 6175 25875 6179 25909
rect 6179 25875 6209 25909
rect 6247 25875 6281 25909
rect 6319 25875 6349 25909
rect 6349 25875 6353 25909
rect 6391 25875 6417 25909
rect 6417 25875 6425 25909
rect 6463 25875 6485 25909
rect 6485 25875 6497 25909
rect 6535 25875 6553 25909
rect 6553 25875 6569 25909
rect 6607 25875 6621 25909
rect 6621 25875 6641 25909
rect 6679 25875 6689 25909
rect 6689 25875 6713 25909
rect 6751 25875 6757 25909
rect 6757 25875 6785 25909
rect 6823 25875 6825 25909
rect 6825 25875 6857 25909
rect 6895 25875 6927 25909
rect 6927 25875 6929 25909
rect 6967 25875 6995 25909
rect 6995 25875 7001 25909
rect 7039 25875 7063 25909
rect 7063 25875 7073 25909
rect 7111 25875 7131 25909
rect 7131 25875 7145 25909
rect 7183 25875 7199 25909
rect 7199 25875 7217 25909
rect 7255 25875 7267 25909
rect 7267 25875 7289 25909
rect 7327 25875 7335 25909
rect 7335 25875 7361 25909
rect 7399 25875 7403 25909
rect 7403 25875 7433 25909
rect 7471 25875 7505 25909
rect 7543 25875 7573 25909
rect 7573 25875 7577 25909
rect 7615 25875 7641 25909
rect 7641 25875 7649 25909
rect 7687 25875 7709 25909
rect 7709 25875 7721 25909
rect 7759 25875 7777 25909
rect 7777 25875 7793 25909
rect 7831 25875 7845 25909
rect 7845 25875 7865 25909
rect 7903 25875 7913 25909
rect 7913 25875 7937 25909
rect 7975 25875 7981 25909
rect 7981 25875 8009 25909
rect 8047 25875 8049 25909
rect 8049 25875 8081 25909
rect 8119 25875 8151 25909
rect 8151 25875 8153 25909
rect 8191 25875 8219 25909
rect 8219 25875 8225 25909
rect 8263 25875 8287 25909
rect 8287 25875 8297 25909
rect 8335 25875 8355 25909
rect 8355 25875 8369 25909
rect 8407 25875 8423 25909
rect 8423 25875 8441 25909
rect 8479 25875 8491 25909
rect 8491 25875 8513 25909
rect 8551 25875 8559 25909
rect 8559 25875 8585 25909
rect 8623 25875 8627 25909
rect 8627 25875 8657 25909
rect 8695 25875 8729 25909
rect 8767 25875 8797 25909
rect 8797 25875 8801 25909
rect 8839 25875 8865 25909
rect 8865 25875 8873 25909
rect 8911 25875 8933 25909
rect 8933 25875 8945 25909
rect 8983 25875 9001 25909
rect 9001 25875 9017 25909
rect 9055 25875 9069 25909
rect 9069 25875 9089 25909
rect 9127 25875 9137 25909
rect 9137 25875 9161 25909
rect 9199 25875 9205 25909
rect 9205 25875 9233 25909
rect 9271 25875 9273 25909
rect 9273 25875 9305 25909
rect 9343 25875 9375 25909
rect 9375 25875 9377 25909
rect 9415 25875 9443 25909
rect 9443 25875 9449 25909
rect 9487 25875 9511 25909
rect 9511 25875 9521 25909
rect 9559 25875 9579 25909
rect 9579 25875 9593 25909
rect 9631 25875 9647 25909
rect 9647 25875 9665 25909
rect 9703 25875 9715 25909
rect 9715 25875 9737 25909
rect 9775 25875 9783 25909
rect 9783 25875 9809 25909
rect 9847 25875 9851 25909
rect 9851 25875 9881 25909
rect 9919 25875 9953 25909
rect 9991 25875 10021 25909
rect 10021 25875 10025 25909
rect 10063 25875 10089 25909
rect 10089 25875 10097 25909
rect 10135 25875 10157 25909
rect 10157 25875 10169 25909
rect 10207 25875 10225 25909
rect 10225 25875 10241 25909
rect 10279 25875 10293 25909
rect 10293 25875 10313 25909
rect 10351 25875 10361 25909
rect 10361 25875 10385 25909
rect 10423 25875 10429 25909
rect 10429 25875 10457 25909
rect 10495 25875 10497 25909
rect 10497 25875 10529 25909
rect 10567 25875 10599 25909
rect 10599 25875 10601 25909
rect 10639 25875 10667 25909
rect 10667 25875 10673 25909
rect 10711 25875 10735 25909
rect 10735 25875 10745 25909
rect 10783 25875 10803 25909
rect 10803 25875 10817 25909
rect 10855 25875 10871 25909
rect 10871 25875 10889 25909
rect 10927 25875 10939 25909
rect 10939 25875 10961 25909
rect 10999 25875 11007 25909
rect 11007 25875 11033 25909
rect 11071 25875 11075 25909
rect 11075 25875 11105 25909
rect 11143 25875 11177 25909
rect 11215 25875 11245 25909
rect 11245 25875 11249 25909
rect 11287 25875 11313 25909
rect 11313 25875 11321 25909
rect 11359 25875 11381 25909
rect 11381 25875 11393 25909
rect 11431 25875 11449 25909
rect 11449 25875 11465 25909
rect 11503 25875 11517 25909
rect 11517 25875 11537 25909
rect 11575 25875 11585 25909
rect 11585 25875 11609 25909
rect 11647 25875 11653 25909
rect 11653 25875 11681 25909
rect 11719 25875 11721 25909
rect 11721 25875 11753 25909
rect 11791 25875 11823 25909
rect 11823 25875 11825 25909
rect 11863 25875 11891 25909
rect 11891 25875 11897 25909
rect 11935 25875 11959 25909
rect 11959 25875 11969 25909
rect 12007 25875 12027 25909
rect 12027 25875 12041 25909
rect 12079 25875 12095 25909
rect 12095 25875 12113 25909
rect 12151 25875 12163 25909
rect 12163 25875 12185 25909
rect 12223 25875 12231 25909
rect 12231 25875 12257 25909
rect 12295 25875 12299 25909
rect 12299 25875 12329 25909
rect 12367 25875 12401 25909
rect 12439 25875 12469 25909
rect 12469 25875 12473 25909
rect 2386 25792 2420 25796
rect 2386 25762 2420 25792
rect 2386 25690 2420 25724
rect 2386 25622 2420 25652
rect 2386 25618 2420 25622
rect 2503 25654 2507 25760
rect 2507 25654 12469 25760
rect 12469 25654 12473 25760
rect 12556 25792 12590 25796
rect 12556 25762 12590 25792
rect 12556 25690 12590 25724
rect 12556 25622 12590 25652
rect 12556 25618 12590 25622
rect 2503 25505 2507 25539
rect 2507 25505 2537 25539
rect 2575 25505 2609 25539
rect 2647 25505 2677 25539
rect 2677 25505 2681 25539
rect 2719 25505 2745 25539
rect 2745 25505 2753 25539
rect 2791 25505 2813 25539
rect 2813 25505 2825 25539
rect 2863 25505 2881 25539
rect 2881 25505 2897 25539
rect 2935 25505 2949 25539
rect 2949 25505 2969 25539
rect 3007 25505 3017 25539
rect 3017 25505 3041 25539
rect 3079 25505 3085 25539
rect 3085 25505 3113 25539
rect 3151 25505 3153 25539
rect 3153 25505 3185 25539
rect 3223 25505 3255 25539
rect 3255 25505 3257 25539
rect 3295 25505 3323 25539
rect 3323 25505 3329 25539
rect 3367 25505 3391 25539
rect 3391 25505 3401 25539
rect 3439 25505 3459 25539
rect 3459 25505 3473 25539
rect 3511 25505 3527 25539
rect 3527 25505 3545 25539
rect 3583 25505 3595 25539
rect 3595 25505 3617 25539
rect 3655 25505 3663 25539
rect 3663 25505 3689 25539
rect 3727 25505 3731 25539
rect 3731 25505 3761 25539
rect 3799 25505 3833 25539
rect 3871 25505 3901 25539
rect 3901 25505 3905 25539
rect 3943 25505 3969 25539
rect 3969 25505 3977 25539
rect 4015 25505 4037 25539
rect 4037 25505 4049 25539
rect 4087 25505 4105 25539
rect 4105 25505 4121 25539
rect 4159 25505 4173 25539
rect 4173 25505 4193 25539
rect 4231 25505 4241 25539
rect 4241 25505 4265 25539
rect 4303 25505 4309 25539
rect 4309 25505 4337 25539
rect 4375 25505 4377 25539
rect 4377 25505 4409 25539
rect 4447 25505 4479 25539
rect 4479 25505 4481 25539
rect 4519 25505 4547 25539
rect 4547 25505 4553 25539
rect 4591 25505 4615 25539
rect 4615 25505 4625 25539
rect 4663 25505 4683 25539
rect 4683 25505 4697 25539
rect 4735 25505 4751 25539
rect 4751 25505 4769 25539
rect 4807 25505 4819 25539
rect 4819 25505 4841 25539
rect 4879 25505 4887 25539
rect 4887 25505 4913 25539
rect 4951 25505 4955 25539
rect 4955 25505 4985 25539
rect 5023 25505 5057 25539
rect 5095 25505 5125 25539
rect 5125 25505 5129 25539
rect 5167 25505 5193 25539
rect 5193 25505 5201 25539
rect 5239 25505 5261 25539
rect 5261 25505 5273 25539
rect 5311 25505 5329 25539
rect 5329 25505 5345 25539
rect 5383 25505 5397 25539
rect 5397 25505 5417 25539
rect 5455 25505 5465 25539
rect 5465 25505 5489 25539
rect 5527 25505 5533 25539
rect 5533 25505 5561 25539
rect 5599 25505 5601 25539
rect 5601 25505 5633 25539
rect 5671 25505 5703 25539
rect 5703 25505 5705 25539
rect 5743 25505 5771 25539
rect 5771 25505 5777 25539
rect 5815 25505 5839 25539
rect 5839 25505 5849 25539
rect 5887 25505 5907 25539
rect 5907 25505 5921 25539
rect 5959 25505 5975 25539
rect 5975 25505 5993 25539
rect 6031 25505 6043 25539
rect 6043 25505 6065 25539
rect 6103 25505 6111 25539
rect 6111 25505 6137 25539
rect 6175 25505 6179 25539
rect 6179 25505 6209 25539
rect 6247 25505 6281 25539
rect 6319 25505 6349 25539
rect 6349 25505 6353 25539
rect 6391 25505 6417 25539
rect 6417 25505 6425 25539
rect 6463 25505 6485 25539
rect 6485 25505 6497 25539
rect 6535 25505 6553 25539
rect 6553 25505 6569 25539
rect 6607 25505 6621 25539
rect 6621 25505 6641 25539
rect 6679 25505 6689 25539
rect 6689 25505 6713 25539
rect 6751 25505 6757 25539
rect 6757 25505 6785 25539
rect 6823 25505 6825 25539
rect 6825 25505 6857 25539
rect 6895 25505 6927 25539
rect 6927 25505 6929 25539
rect 6967 25505 6995 25539
rect 6995 25505 7001 25539
rect 7039 25505 7063 25539
rect 7063 25505 7073 25539
rect 7111 25505 7131 25539
rect 7131 25505 7145 25539
rect 7183 25505 7199 25539
rect 7199 25505 7217 25539
rect 7255 25505 7267 25539
rect 7267 25505 7289 25539
rect 7327 25505 7335 25539
rect 7335 25505 7361 25539
rect 7399 25505 7403 25539
rect 7403 25505 7433 25539
rect 7471 25505 7505 25539
rect 7543 25505 7573 25539
rect 7573 25505 7577 25539
rect 7615 25505 7641 25539
rect 7641 25505 7649 25539
rect 7687 25505 7709 25539
rect 7709 25505 7721 25539
rect 7759 25505 7777 25539
rect 7777 25505 7793 25539
rect 7831 25505 7845 25539
rect 7845 25505 7865 25539
rect 7903 25505 7913 25539
rect 7913 25505 7937 25539
rect 7975 25505 7981 25539
rect 7981 25505 8009 25539
rect 8047 25505 8049 25539
rect 8049 25505 8081 25539
rect 8119 25505 8151 25539
rect 8151 25505 8153 25539
rect 8191 25505 8219 25539
rect 8219 25505 8225 25539
rect 8263 25505 8287 25539
rect 8287 25505 8297 25539
rect 8335 25505 8355 25539
rect 8355 25505 8369 25539
rect 8407 25505 8423 25539
rect 8423 25505 8441 25539
rect 8479 25505 8491 25539
rect 8491 25505 8513 25539
rect 8551 25505 8559 25539
rect 8559 25505 8585 25539
rect 8623 25505 8627 25539
rect 8627 25505 8657 25539
rect 8695 25505 8729 25539
rect 8767 25505 8797 25539
rect 8797 25505 8801 25539
rect 8839 25505 8865 25539
rect 8865 25505 8873 25539
rect 8911 25505 8933 25539
rect 8933 25505 8945 25539
rect 8983 25505 9001 25539
rect 9001 25505 9017 25539
rect 9055 25505 9069 25539
rect 9069 25505 9089 25539
rect 9127 25505 9137 25539
rect 9137 25505 9161 25539
rect 9199 25505 9205 25539
rect 9205 25505 9233 25539
rect 9271 25505 9273 25539
rect 9273 25505 9305 25539
rect 9343 25505 9375 25539
rect 9375 25505 9377 25539
rect 9415 25505 9443 25539
rect 9443 25505 9449 25539
rect 9487 25505 9511 25539
rect 9511 25505 9521 25539
rect 9559 25505 9579 25539
rect 9579 25505 9593 25539
rect 9631 25505 9647 25539
rect 9647 25505 9665 25539
rect 9703 25505 9715 25539
rect 9715 25505 9737 25539
rect 9775 25505 9783 25539
rect 9783 25505 9809 25539
rect 9847 25505 9851 25539
rect 9851 25505 9881 25539
rect 9919 25505 9953 25539
rect 9991 25505 10021 25539
rect 10021 25505 10025 25539
rect 10063 25505 10089 25539
rect 10089 25505 10097 25539
rect 10135 25505 10157 25539
rect 10157 25505 10169 25539
rect 10207 25505 10225 25539
rect 10225 25505 10241 25539
rect 10279 25505 10293 25539
rect 10293 25505 10313 25539
rect 10351 25505 10361 25539
rect 10361 25505 10385 25539
rect 10423 25505 10429 25539
rect 10429 25505 10457 25539
rect 10495 25505 10497 25539
rect 10497 25505 10529 25539
rect 10567 25505 10599 25539
rect 10599 25505 10601 25539
rect 10639 25505 10667 25539
rect 10667 25505 10673 25539
rect 10711 25505 10735 25539
rect 10735 25505 10745 25539
rect 10783 25505 10803 25539
rect 10803 25505 10817 25539
rect 10855 25505 10871 25539
rect 10871 25505 10889 25539
rect 10927 25505 10939 25539
rect 10939 25505 10961 25539
rect 10999 25505 11007 25539
rect 11007 25505 11033 25539
rect 11071 25505 11075 25539
rect 11075 25505 11105 25539
rect 11143 25505 11177 25539
rect 11215 25505 11245 25539
rect 11245 25505 11249 25539
rect 11287 25505 11313 25539
rect 11313 25505 11321 25539
rect 11359 25505 11381 25539
rect 11381 25505 11393 25539
rect 11431 25505 11449 25539
rect 11449 25505 11465 25539
rect 11503 25505 11517 25539
rect 11517 25505 11537 25539
rect 11575 25505 11585 25539
rect 11585 25505 11609 25539
rect 11647 25505 11653 25539
rect 11653 25505 11681 25539
rect 11719 25505 11721 25539
rect 11721 25505 11753 25539
rect 11791 25505 11823 25539
rect 11823 25505 11825 25539
rect 11863 25505 11891 25539
rect 11891 25505 11897 25539
rect 11935 25505 11959 25539
rect 11959 25505 11969 25539
rect 12007 25505 12027 25539
rect 12027 25505 12041 25539
rect 12079 25505 12095 25539
rect 12095 25505 12113 25539
rect 12151 25505 12163 25539
rect 12163 25505 12185 25539
rect 12223 25505 12231 25539
rect 12231 25505 12257 25539
rect 12295 25505 12299 25539
rect 12299 25505 12329 25539
rect 12367 25505 12401 25539
rect 12439 25505 12469 25539
rect 12469 25505 12473 25539
rect 12834 26067 13228 26087
rect 12834 25353 12844 26067
rect 12844 25353 13218 26067
rect 13218 25353 13228 26067
rect 12834 25333 13228 25353
rect 2251 25219 12725 25229
rect 2251 24845 2269 25219
rect 2269 24845 12707 25219
rect 12707 24845 12725 25219
rect 2251 24835 12725 24845
rect 1153 24751 1187 24775
rect 1153 24741 1187 24751
rect 1153 24683 1187 24703
rect 1153 24669 1187 24683
rect 1153 24615 1187 24631
rect 1153 24597 1187 24615
rect 1153 24547 1187 24559
rect 1153 24525 1187 24547
rect 1153 24479 1187 24487
rect 1153 24453 1187 24479
rect 1153 24411 1187 24415
rect 1153 24381 1187 24411
rect 1153 24309 1187 24343
rect 1153 24241 1187 24271
rect 1153 24237 1187 24241
rect 1153 24173 1187 24199
rect 1153 24165 1187 24173
rect 1153 24105 1187 24127
rect 1153 24093 1187 24105
rect 1153 24037 1187 24055
rect 1153 24021 1187 24037
rect 1153 23969 1187 23983
rect 1153 23949 1187 23969
rect 1153 23901 1187 23911
rect 1153 23877 1187 23901
rect 1153 23833 1187 23839
rect 1153 23805 1187 23833
rect 1153 23765 1187 23767
rect 1153 23733 1187 23765
rect 1153 23663 1187 23695
rect 1153 23661 1187 23663
rect 1153 23595 1187 23623
rect 1153 23589 1187 23595
rect 1153 23527 1187 23551
rect 1153 23517 1187 23527
rect 1153 23459 1187 23479
rect 1153 23445 1187 23459
rect 1153 23391 1187 23407
rect 1153 23373 1187 23391
rect 1153 23323 1187 23335
rect 1153 23301 1187 23323
rect 1153 23255 1187 23263
rect 1153 23229 1187 23255
rect 1153 23187 1187 23191
rect 1153 23157 1187 23187
rect 1153 23085 1187 23119
rect 1153 23017 1187 23047
rect 1153 23013 1187 23017
rect 1153 22949 1187 22975
rect 1153 22941 1187 22949
rect 1153 22881 1187 22903
rect 1153 22869 1187 22881
rect 1153 22813 1187 22831
rect 1153 22797 1187 22813
rect 1153 22745 1187 22759
rect 1153 22725 1187 22745
rect 1153 22677 1187 22687
rect 1153 22653 1187 22677
rect 1153 22609 1187 22615
rect 1153 22581 1187 22609
rect 1153 22541 1187 22543
rect 1153 22509 1187 22541
rect 1153 22439 1187 22471
rect 1153 22437 1187 22439
rect 1153 22371 1187 22399
rect 1153 22365 1187 22371
rect 1153 22303 1187 22327
rect 1153 22293 1187 22303
rect 1153 22235 1187 22255
rect 1153 22221 1187 22235
rect 1153 22167 1187 22183
rect 1153 22149 1187 22167
rect 1153 22099 1187 22111
rect 1153 22077 1187 22099
rect 1153 22031 1187 22039
rect 1153 22005 1187 22031
rect 1153 21963 1187 21967
rect 1153 21933 1187 21963
rect 1153 21861 1187 21895
rect 1153 21793 1187 21823
rect 1153 21789 1187 21793
rect 1153 21725 1187 21751
rect 1153 21717 1187 21725
rect 1153 21657 1187 21679
rect 1153 21645 1187 21657
rect 1153 21589 1187 21607
rect 1153 21573 1187 21589
rect 1153 21521 1187 21535
rect 1153 21501 1187 21521
rect 1153 21453 1187 21463
rect 1153 21429 1187 21453
rect 1153 21385 1187 21391
rect 1153 21357 1187 21385
rect 1153 21317 1187 21319
rect 1153 21285 1187 21317
rect 1153 21215 1187 21247
rect 1153 21213 1187 21215
rect 1153 21147 1187 21175
rect 1153 21141 1187 21147
rect 1153 21079 1187 21103
rect 1153 21069 1187 21079
rect 1153 21011 1187 21031
rect 1153 20997 1187 21011
rect 1153 20943 1187 20959
rect 1153 20925 1187 20943
rect 1153 20875 1187 20887
rect 1153 20853 1187 20875
rect 1153 20807 1187 20815
rect 1153 20781 1187 20807
rect 1153 20739 1187 20743
rect 1153 20709 1187 20739
rect 1153 20637 1187 20671
rect 1153 20569 1187 20599
rect 1153 20565 1187 20569
rect 1153 20501 1187 20527
rect 1153 20493 1187 20501
rect 1153 20433 1187 20455
rect 1153 20421 1187 20433
rect 1153 20365 1187 20383
rect 1153 20349 1187 20365
rect 1153 20297 1187 20311
rect 1153 20277 1187 20297
rect 1153 20229 1187 20239
rect 1153 20205 1187 20229
rect 1153 20161 1187 20167
rect 1153 20133 1187 20161
rect 1153 20093 1187 20095
rect 1153 20061 1187 20093
rect 1153 19991 1187 20023
rect 1153 19989 1187 19991
rect 1153 19923 1187 19951
rect 1153 19917 1187 19923
rect 1153 19855 1187 19879
rect 1153 19845 1187 19855
rect 1153 19787 1187 19807
rect 1153 19773 1187 19787
rect 1153 19719 1187 19735
rect 1153 19701 1187 19719
rect 1153 19651 1187 19663
rect 1153 19629 1187 19651
rect 1153 19583 1187 19591
rect 1153 19557 1187 19583
rect 1153 19515 1187 19519
rect 1153 19485 1187 19515
rect 1153 19413 1187 19447
rect 1153 19345 1187 19375
rect 1153 19341 1187 19345
rect 1153 19277 1187 19303
rect 1153 19269 1187 19277
rect 1153 19209 1187 19231
rect 1153 19197 1187 19209
rect 1153 19141 1187 19159
rect 1153 19125 1187 19141
rect 1153 19073 1187 19087
rect 1153 19053 1187 19073
rect 1153 19005 1187 19015
rect 1153 18981 1187 19005
rect 1153 18937 1187 18943
rect 1153 18909 1187 18937
rect 1153 18869 1187 18871
rect 1153 18837 1187 18869
rect 1153 18767 1187 18799
rect 1153 18765 1187 18767
rect 1153 18699 1187 18727
rect 1153 18693 1187 18699
rect 1153 18631 1187 18655
rect 1153 18621 1187 18631
rect 1153 18563 1187 18583
rect 1153 18549 1187 18563
rect 1153 18495 1187 18511
rect 1153 18477 1187 18495
rect 1153 18427 1187 18439
rect 1153 18405 1187 18427
rect 1153 18359 1187 18367
rect 1153 18333 1187 18359
rect 1153 18291 1187 18295
rect 1153 18261 1187 18291
rect 1153 18189 1187 18223
rect 1153 18121 1187 18151
rect 1153 18117 1187 18121
rect 1153 18053 1187 18079
rect 1153 18045 1187 18053
rect 1153 17985 1187 18007
rect 1153 17973 1187 17985
rect 1153 17917 1187 17935
rect 1153 17901 1187 17917
rect 1153 17849 1187 17863
rect 1153 17829 1187 17849
rect 1153 17781 1187 17791
rect 1153 17757 1187 17781
rect 1153 17713 1187 17719
rect 1153 17685 1187 17713
rect 1153 17645 1187 17647
rect 1153 17613 1187 17645
rect 1153 17543 1187 17575
rect 1153 17541 1187 17543
rect 1153 17475 1187 17503
rect 1153 17469 1187 17475
rect 1153 17407 1187 17431
rect 1153 17397 1187 17407
rect 1153 17339 1187 17359
rect 1153 17325 1187 17339
rect 1153 17271 1187 17287
rect 1153 17253 1187 17271
rect 1153 17203 1187 17215
rect 1153 17181 1187 17203
rect 1153 17135 1187 17143
rect 1153 17109 1187 17135
rect 1153 17067 1187 17071
rect 1153 17037 1187 17067
rect 1153 16965 1187 16999
rect 1153 16897 1187 16927
rect 1153 16893 1187 16897
rect 1153 16829 1187 16855
rect 1153 16821 1187 16829
rect 1153 16761 1187 16783
rect 1153 16749 1187 16761
rect 1153 16693 1187 16711
rect 1153 16677 1187 16693
rect 1153 16625 1187 16639
rect 1153 16605 1187 16625
rect 1153 16557 1187 16567
rect 1153 16533 1187 16557
rect 1153 16489 1187 16495
rect 1153 16461 1187 16489
rect 1153 16421 1187 16423
rect 1153 16389 1187 16421
rect 1153 16319 1187 16351
rect 1153 16317 1187 16319
rect 1153 16251 1187 16279
rect 1153 16245 1187 16251
rect 1153 16183 1187 16207
rect 1153 16173 1187 16183
rect 1153 16115 1187 16135
rect 1153 16101 1187 16115
rect 1153 16047 1187 16063
rect 1153 16029 1187 16047
rect 1153 15979 1187 15991
rect 1153 15957 1187 15979
rect 1153 15911 1187 15919
rect 1153 15885 1187 15911
rect 1153 15843 1187 15847
rect 1153 15813 1187 15843
rect 1153 15741 1187 15775
rect 1153 15673 1187 15703
rect 1153 15669 1187 15673
rect 1153 15605 1187 15631
rect 1153 15597 1187 15605
rect 1153 15537 1187 15559
rect 1153 15525 1187 15537
rect 1153 15469 1187 15487
rect 1153 15453 1187 15469
rect 1153 15401 1187 15415
rect 1153 15381 1187 15401
rect 13801 23386 13835 23410
rect 13801 23376 13835 23386
rect 13801 23318 13835 23338
rect 13801 23304 13835 23318
rect 13801 23250 13835 23266
rect 13801 23232 13835 23250
rect 13801 23182 13835 23194
rect 13801 23160 13835 23182
rect 13801 23114 13835 23122
rect 13801 23088 13835 23114
rect 13801 23046 13835 23050
rect 13801 23016 13835 23046
rect 13801 22944 13835 22978
rect 13801 22876 13835 22906
rect 13801 22872 13835 22876
rect 13801 22808 13835 22834
rect 13801 22800 13835 22808
rect 13801 22740 13835 22762
rect 13801 22728 13835 22740
rect 13801 22672 13835 22690
rect 13801 22656 13835 22672
rect 13801 22604 13835 22618
rect 13801 22584 13835 22604
rect 13801 22536 13835 22546
rect 13801 22512 13835 22536
rect 13801 22468 13835 22474
rect 13801 22440 13835 22468
rect 13801 22400 13835 22402
rect 13801 22368 13835 22400
rect 13801 22298 13835 22330
rect 13801 22296 13835 22298
rect 13801 22230 13835 22258
rect 13801 22224 13835 22230
rect 13801 22162 13835 22186
rect 13801 22152 13835 22162
rect 13801 22094 13835 22114
rect 13801 22080 13835 22094
rect 13801 22026 13835 22042
rect 13801 22008 13835 22026
rect 13801 21958 13835 21970
rect 13801 21936 13835 21958
rect 13801 21890 13835 21898
rect 13801 21864 13835 21890
rect 13801 21822 13835 21826
rect 13801 21792 13835 21822
rect 13801 21720 13835 21754
rect 13801 21652 13835 21682
rect 13801 21648 13835 21652
rect 13801 21584 13835 21610
rect 13801 21576 13835 21584
rect 13801 21516 13835 21538
rect 13801 21504 13835 21516
rect 13801 21448 13835 21466
rect 13801 21432 13835 21448
rect 13801 21380 13835 21394
rect 13801 21360 13835 21380
rect 13801 21312 13835 21322
rect 13801 21288 13835 21312
rect 13801 21244 13835 21250
rect 13801 21216 13835 21244
rect 13801 21176 13835 21178
rect 13801 21144 13835 21176
rect 13801 21074 13835 21106
rect 13801 21072 13835 21074
rect 13801 21006 13835 21034
rect 13801 21000 13835 21006
rect 13801 20938 13835 20962
rect 13801 20928 13835 20938
rect 13801 20870 13835 20890
rect 13801 20856 13835 20870
rect 13801 20802 13835 20818
rect 13801 20784 13835 20802
rect 13801 20734 13835 20746
rect 13801 20712 13835 20734
rect 13801 20666 13835 20674
rect 13801 20640 13835 20666
rect 13801 20598 13835 20602
rect 13801 20568 13835 20598
rect 13801 20496 13835 20530
rect 13801 20428 13835 20458
rect 13801 20424 13835 20428
rect 13801 20360 13835 20386
rect 13801 20352 13835 20360
rect 13801 20292 13835 20314
rect 13801 20280 13835 20292
rect 13801 20224 13835 20242
rect 13801 20208 13835 20224
rect 13801 20156 13835 20170
rect 13801 20136 13835 20156
rect 13801 20088 13835 20098
rect 13801 20064 13835 20088
rect 13801 20020 13835 20026
rect 13801 19992 13835 20020
rect 13801 19952 13835 19954
rect 13801 19920 13835 19952
rect 13801 19850 13835 19882
rect 13801 19848 13835 19850
rect 13801 19782 13835 19810
rect 13801 19776 13835 19782
rect 13801 19714 13835 19738
rect 13801 19704 13835 19714
rect 13801 19646 13835 19666
rect 13801 19632 13835 19646
rect 13801 19578 13835 19594
rect 13801 19560 13835 19578
rect 13801 19510 13835 19522
rect 13801 19488 13835 19510
rect 13801 19442 13835 19450
rect 13801 19416 13835 19442
rect 13801 19374 13835 19378
rect 13801 19344 13835 19374
rect 13801 19272 13835 19306
rect 13801 19204 13835 19234
rect 13801 19200 13835 19204
rect 13801 19136 13835 19162
rect 13801 19128 13835 19136
rect 13801 19068 13835 19090
rect 13801 19056 13835 19068
rect 13801 19000 13835 19018
rect 13801 18984 13835 19000
rect 13801 18932 13835 18946
rect 13801 18912 13835 18932
rect 13801 18864 13835 18874
rect 13801 18840 13835 18864
rect 13801 18796 13835 18802
rect 13801 18768 13835 18796
rect 13801 18728 13835 18730
rect 13801 18696 13835 18728
rect 13801 18626 13835 18658
rect 13801 18624 13835 18626
rect 13801 18558 13835 18586
rect 13801 18552 13835 18558
rect 13801 18490 13835 18514
rect 13801 18480 13835 18490
rect 13801 18422 13835 18442
rect 13801 18408 13835 18422
rect 13801 18354 13835 18370
rect 13801 18336 13835 18354
rect 13801 18286 13835 18298
rect 13801 18264 13835 18286
rect 13801 18218 13835 18226
rect 13801 18192 13835 18218
rect 13801 18150 13835 18154
rect 13801 18120 13835 18150
rect 13801 18048 13835 18082
rect 13801 17980 13835 18010
rect 13801 17976 13835 17980
rect 13801 17912 13835 17938
rect 13801 17904 13835 17912
rect 13801 17844 13835 17866
rect 13801 17832 13835 17844
rect 13801 17776 13835 17794
rect 13801 17760 13835 17776
rect 13801 17708 13835 17722
rect 13801 17688 13835 17708
rect 13801 17640 13835 17650
rect 13801 17616 13835 17640
rect 13801 17572 13835 17578
rect 13801 17544 13835 17572
rect 13801 17504 13835 17506
rect 13801 17472 13835 17504
rect 13801 17402 13835 17434
rect 13801 17400 13835 17402
rect 13801 17334 13835 17362
rect 13801 17328 13835 17334
rect 13801 17266 13835 17290
rect 13801 17256 13835 17266
rect 13801 17198 13835 17218
rect 13801 17184 13835 17198
rect 13801 17130 13835 17146
rect 13801 17112 13835 17130
rect 13801 17062 13835 17074
rect 13801 17040 13835 17062
rect 13801 16994 13835 17002
rect 13801 16968 13835 16994
rect 13801 16926 13835 16930
rect 13801 16896 13835 16926
rect 13801 16824 13835 16858
rect 13801 16756 13835 16786
rect 13801 16752 13835 16756
rect 13801 16688 13835 16714
rect 13801 16680 13835 16688
rect 13801 16620 13835 16642
rect 13801 16608 13835 16620
rect 13801 16552 13835 16570
rect 13801 16536 13835 16552
rect 13801 16484 13835 16498
rect 13801 16464 13835 16484
rect 13801 16416 13835 16426
rect 13801 16392 13835 16416
rect 13801 16348 13835 16354
rect 13801 16320 13835 16348
rect 13801 16280 13835 16282
rect 13801 16248 13835 16280
rect 13801 16178 13835 16210
rect 13801 16176 13835 16178
rect 13801 16110 13835 16138
rect 13801 16104 13835 16110
rect 13801 16042 13835 16066
rect 13801 16032 13835 16042
rect 13801 15974 13835 15994
rect 13801 15960 13835 15974
rect 13801 15906 13835 15922
rect 13801 15888 13835 15906
rect 13801 15838 13835 15850
rect 13801 15816 13835 15838
rect 13801 15770 13835 15778
rect 13801 15744 13835 15770
rect 13801 15702 13835 15706
rect 13801 15672 13835 15702
rect 13801 15600 13835 15634
rect 13801 15532 13835 15562
rect 13801 15528 13835 15532
rect 13801 15464 13835 15490
rect 13801 15456 13835 15464
rect 13801 15396 13835 15418
rect 13801 15384 13835 15396
rect 1290 15257 1294 15291
rect 1294 15257 1324 15291
rect 1362 15257 1396 15291
rect 1434 15257 1464 15291
rect 1464 15257 1468 15291
rect 1506 15257 1532 15291
rect 1532 15257 1540 15291
rect 1578 15257 1600 15291
rect 1600 15257 1612 15291
rect 1650 15257 1668 15291
rect 1668 15257 1684 15291
rect 1722 15257 1736 15291
rect 1736 15257 1756 15291
rect 1794 15257 1804 15291
rect 1804 15257 1828 15291
rect 1866 15257 1872 15291
rect 1872 15257 1900 15291
rect 1938 15257 1940 15291
rect 1940 15257 1972 15291
rect 2010 15257 2042 15291
rect 2042 15257 2044 15291
rect 2082 15257 2110 15291
rect 2110 15257 2116 15291
rect 2154 15257 2178 15291
rect 2178 15257 2188 15291
rect 2226 15257 2246 15291
rect 2246 15257 2260 15291
rect 2298 15257 2314 15291
rect 2314 15257 2332 15291
rect 2370 15257 2382 15291
rect 2382 15257 2404 15291
rect 2442 15257 2450 15291
rect 2450 15257 2476 15291
rect 2514 15257 2518 15291
rect 2518 15257 2548 15291
rect 2586 15257 2620 15291
rect 2658 15257 2688 15291
rect 2688 15257 2692 15291
rect 2730 15257 2756 15291
rect 2756 15257 2764 15291
rect 2802 15257 2824 15291
rect 2824 15257 2836 15291
rect 2874 15257 2892 15291
rect 2892 15257 2908 15291
rect 2946 15257 2960 15291
rect 2960 15257 2980 15291
rect 3018 15257 3028 15291
rect 3028 15257 3052 15291
rect 3090 15257 3096 15291
rect 3096 15257 3124 15291
rect 3162 15257 3164 15291
rect 3164 15257 3196 15291
rect 3234 15257 3266 15291
rect 3266 15257 3268 15291
rect 3306 15257 3334 15291
rect 3334 15257 3340 15291
rect 3378 15257 3402 15291
rect 3402 15257 3412 15291
rect 3450 15257 3470 15291
rect 3470 15257 3484 15291
rect 3522 15257 3538 15291
rect 3538 15257 3556 15291
rect 3594 15257 3606 15291
rect 3606 15257 3628 15291
rect 3666 15257 3674 15291
rect 3674 15257 3700 15291
rect 3738 15257 3742 15291
rect 3742 15257 3772 15291
rect 3810 15257 3844 15291
rect 3882 15257 3912 15291
rect 3912 15257 3916 15291
rect 3954 15257 3980 15291
rect 3980 15257 3988 15291
rect 4026 15257 4048 15291
rect 4048 15257 4060 15291
rect 4098 15257 4116 15291
rect 4116 15257 4132 15291
rect 4170 15257 4184 15291
rect 4184 15257 4204 15291
rect 4242 15257 4252 15291
rect 4252 15257 4276 15291
rect 4314 15257 4320 15291
rect 4320 15257 4348 15291
rect 4386 15257 4388 15291
rect 4388 15257 4420 15291
rect 4458 15257 4490 15291
rect 4490 15257 4492 15291
rect 4530 15257 4558 15291
rect 4558 15257 4564 15291
rect 4602 15257 4626 15291
rect 4626 15257 4636 15291
rect 4674 15257 4694 15291
rect 4694 15257 4708 15291
rect 4746 15257 4762 15291
rect 4762 15257 4780 15291
rect 4818 15257 4830 15291
rect 4830 15257 4852 15291
rect 4890 15257 4898 15291
rect 4898 15257 4924 15291
rect 4962 15257 4966 15291
rect 4966 15257 4996 15291
rect 5034 15257 5068 15291
rect 5106 15257 5136 15291
rect 5136 15257 5140 15291
rect 5178 15257 5204 15291
rect 5204 15257 5212 15291
rect 5250 15257 5272 15291
rect 5272 15257 5284 15291
rect 5322 15257 5340 15291
rect 5340 15257 5356 15291
rect 5394 15257 5408 15291
rect 5408 15257 5428 15291
rect 5466 15257 5476 15291
rect 5476 15257 5500 15291
rect 5538 15257 5544 15291
rect 5544 15257 5572 15291
rect 5610 15257 5612 15291
rect 5612 15257 5644 15291
rect 5682 15257 5714 15291
rect 5714 15257 5716 15291
rect 5754 15257 5782 15291
rect 5782 15257 5788 15291
rect 5826 15257 5850 15291
rect 5850 15257 5860 15291
rect 5898 15257 5918 15291
rect 5918 15257 5932 15291
rect 5970 15257 5986 15291
rect 5986 15257 6004 15291
rect 6042 15257 6054 15291
rect 6054 15257 6076 15291
rect 6114 15257 6122 15291
rect 6122 15257 6148 15291
rect 6186 15257 6190 15291
rect 6190 15257 6220 15291
rect 6258 15257 6292 15291
rect 6330 15257 6360 15291
rect 6360 15257 6364 15291
rect 6402 15257 6428 15291
rect 6428 15257 6436 15291
rect 6474 15257 6496 15291
rect 6496 15257 6508 15291
rect 6546 15257 6564 15291
rect 6564 15257 6580 15291
rect 6618 15257 6632 15291
rect 6632 15257 6652 15291
rect 6690 15257 6700 15291
rect 6700 15257 6724 15291
rect 6762 15257 6768 15291
rect 6768 15257 6796 15291
rect 6834 15257 6836 15291
rect 6836 15257 6868 15291
rect 6906 15257 6938 15291
rect 6938 15257 6940 15291
rect 6978 15257 7006 15291
rect 7006 15257 7012 15291
rect 7050 15257 7074 15291
rect 7074 15257 7084 15291
rect 7122 15257 7142 15291
rect 7142 15257 7156 15291
rect 7194 15257 7210 15291
rect 7210 15257 7228 15291
rect 7266 15257 7278 15291
rect 7278 15257 7300 15291
rect 7338 15257 7346 15291
rect 7346 15257 7372 15291
rect 7410 15257 7414 15291
rect 7414 15257 7444 15291
rect 7482 15257 7516 15291
rect 7554 15257 7584 15291
rect 7584 15257 7588 15291
rect 7626 15257 7652 15291
rect 7652 15257 7660 15291
rect 7698 15257 7720 15291
rect 7720 15257 7732 15291
rect 7770 15257 7788 15291
rect 7788 15257 7804 15291
rect 7842 15257 7856 15291
rect 7856 15257 7876 15291
rect 7914 15257 7924 15291
rect 7924 15257 7948 15291
rect 7986 15257 7992 15291
rect 7992 15257 8020 15291
rect 8058 15257 8060 15291
rect 8060 15257 8092 15291
rect 8130 15257 8162 15291
rect 8162 15257 8164 15291
rect 8202 15257 8230 15291
rect 8230 15257 8236 15291
rect 8274 15257 8298 15291
rect 8298 15257 8308 15291
rect 8346 15257 8366 15291
rect 8366 15257 8380 15291
rect 8418 15257 8434 15291
rect 8434 15257 8452 15291
rect 8490 15257 8502 15291
rect 8502 15257 8524 15291
rect 8562 15257 8570 15291
rect 8570 15257 8596 15291
rect 8634 15257 8638 15291
rect 8638 15257 8668 15291
rect 8706 15257 8740 15291
rect 8778 15257 8808 15291
rect 8808 15257 8812 15291
rect 8850 15257 8876 15291
rect 8876 15257 8884 15291
rect 8922 15257 8944 15291
rect 8944 15257 8956 15291
rect 8994 15257 9012 15291
rect 9012 15257 9028 15291
rect 9066 15257 9080 15291
rect 9080 15257 9100 15291
rect 9138 15257 9148 15291
rect 9148 15257 9172 15291
rect 9210 15257 9216 15291
rect 9216 15257 9244 15291
rect 9282 15257 9284 15291
rect 9284 15257 9316 15291
rect 9354 15257 9386 15291
rect 9386 15257 9388 15291
rect 9426 15257 9454 15291
rect 9454 15257 9460 15291
rect 9498 15257 9522 15291
rect 9522 15257 9532 15291
rect 9570 15257 9590 15291
rect 9590 15257 9604 15291
rect 9642 15257 9658 15291
rect 9658 15257 9676 15291
rect 9714 15257 9726 15291
rect 9726 15257 9748 15291
rect 9786 15257 9794 15291
rect 9794 15257 9820 15291
rect 9858 15257 9862 15291
rect 9862 15257 9892 15291
rect 9930 15257 9964 15291
rect 10002 15257 10032 15291
rect 10032 15257 10036 15291
rect 10074 15257 10100 15291
rect 10100 15257 10108 15291
rect 10146 15257 10168 15291
rect 10168 15257 10180 15291
rect 10218 15257 10236 15291
rect 10236 15257 10252 15291
rect 10290 15257 10304 15291
rect 10304 15257 10324 15291
rect 10362 15257 10372 15291
rect 10372 15257 10396 15291
rect 10434 15257 10440 15291
rect 10440 15257 10468 15291
rect 10506 15257 10508 15291
rect 10508 15257 10540 15291
rect 10578 15257 10610 15291
rect 10610 15257 10612 15291
rect 10650 15257 10678 15291
rect 10678 15257 10684 15291
rect 10722 15257 10746 15291
rect 10746 15257 10756 15291
rect 10794 15257 10814 15291
rect 10814 15257 10828 15291
rect 10866 15257 10882 15291
rect 10882 15257 10900 15291
rect 10938 15257 10950 15291
rect 10950 15257 10972 15291
rect 11010 15257 11018 15291
rect 11018 15257 11044 15291
rect 11082 15257 11086 15291
rect 11086 15257 11116 15291
rect 11154 15257 11188 15291
rect 11226 15257 11256 15291
rect 11256 15257 11260 15291
rect 11298 15257 11324 15291
rect 11324 15257 11332 15291
rect 11370 15257 11392 15291
rect 11392 15257 11404 15291
rect 11442 15257 11460 15291
rect 11460 15257 11476 15291
rect 11514 15257 11528 15291
rect 11528 15257 11548 15291
rect 11586 15257 11596 15291
rect 11596 15257 11620 15291
rect 11658 15257 11664 15291
rect 11664 15257 11692 15291
rect 11730 15257 11732 15291
rect 11732 15257 11764 15291
rect 11802 15257 11834 15291
rect 11834 15257 11836 15291
rect 11874 15257 11902 15291
rect 11902 15257 11908 15291
rect 11946 15257 11970 15291
rect 11970 15257 11980 15291
rect 12018 15257 12038 15291
rect 12038 15257 12052 15291
rect 12090 15257 12106 15291
rect 12106 15257 12124 15291
rect 12162 15257 12174 15291
rect 12174 15257 12196 15291
rect 12234 15257 12242 15291
rect 12242 15257 12268 15291
rect 12306 15257 12310 15291
rect 12310 15257 12340 15291
rect 12378 15257 12412 15291
rect 12450 15257 12480 15291
rect 12480 15257 12484 15291
rect 12522 15257 12548 15291
rect 12548 15257 12556 15291
rect 12594 15257 12616 15291
rect 12616 15257 12628 15291
rect 12666 15257 12684 15291
rect 12684 15257 12700 15291
rect 12738 15257 12752 15291
rect 12752 15257 12772 15291
rect 12810 15257 12820 15291
rect 12820 15257 12844 15291
rect 12882 15257 12888 15291
rect 12888 15257 12916 15291
rect 12954 15257 12956 15291
rect 12956 15257 12988 15291
rect 13026 15257 13058 15291
rect 13058 15257 13060 15291
rect 13098 15257 13126 15291
rect 13126 15257 13132 15291
rect 13170 15257 13194 15291
rect 13194 15257 13204 15291
rect 13242 15257 13262 15291
rect 13262 15257 13276 15291
rect 13314 15257 13330 15291
rect 13330 15257 13348 15291
rect 13386 15257 13398 15291
rect 13398 15257 13420 15291
rect 13458 15257 13466 15291
rect 13466 15257 13492 15291
rect 13530 15257 13534 15291
rect 13534 15257 13564 15291
rect 13602 15257 13636 15291
rect 13674 15257 13704 15291
rect 13704 15257 13708 15291
rect 14114 34720 14148 34754
rect 14114 34648 14148 34682
rect 14114 34576 14148 34610
rect 14114 34504 14148 34538
rect 14114 34432 14148 34466
rect 14114 34360 14148 34394
rect 14114 34288 14148 34322
rect 14114 34216 14148 34250
rect 14114 34144 14148 34178
rect 14114 34072 14148 34106
rect 14114 34000 14148 34034
rect 14114 33928 14148 33962
rect 14114 33856 14148 33890
rect 14114 33784 14148 33818
rect 14114 33712 14148 33746
rect 14114 33640 14148 33674
rect 14114 33568 14148 33602
rect 14114 33496 14148 33530
rect 14114 33424 14148 33458
rect 14114 33352 14148 33386
rect 14114 33280 14148 33314
rect 14114 33208 14148 33242
rect 14114 33136 14148 33170
rect 14114 33064 14148 33098
rect 14114 32992 14148 33026
rect 14114 32920 14148 32954
rect 14114 32848 14148 32882
rect 14114 32776 14148 32810
rect 14114 32704 14148 32738
rect 14114 32632 14148 32666
rect 14114 32560 14148 32594
rect 14114 32488 14148 32522
rect 14114 32416 14148 32450
rect 14114 32344 14148 32378
rect 14114 32272 14148 32306
rect 14114 32200 14148 32234
rect 14114 32128 14148 32162
rect 14114 32056 14148 32090
rect 14114 31984 14148 32018
rect 14114 31912 14148 31946
rect 14114 31840 14148 31874
rect 14114 31768 14148 31802
rect 14114 31696 14148 31730
rect 14114 31624 14148 31658
rect 14114 31552 14148 31586
rect 14114 31480 14148 31514
rect 14114 31408 14148 31442
rect 14114 31336 14148 31370
rect 14114 31264 14148 31298
rect 14114 31192 14148 31226
rect 14114 31120 14148 31154
rect 14114 31048 14148 31082
rect 14114 30976 14148 31010
rect 14114 30904 14148 30938
rect 14114 30832 14148 30866
rect 14114 30760 14148 30794
rect 14114 30688 14148 30722
rect 14114 30616 14148 30650
rect 14114 30544 14148 30578
rect 14114 30472 14148 30506
rect 14114 30400 14148 30434
rect 14114 30328 14148 30362
rect 14114 30256 14148 30290
rect 14114 30184 14148 30218
rect 14114 30112 14148 30146
rect 14114 30040 14148 30074
rect 14114 29968 14148 30002
rect 14114 29896 14148 29930
rect 14114 29824 14148 29858
rect 14114 29752 14148 29786
rect 14114 29680 14148 29714
rect 14114 29608 14148 29642
rect 14114 29536 14148 29570
rect 14114 29464 14148 29498
rect 14114 29392 14148 29426
rect 14114 29320 14148 29354
rect 14114 29248 14148 29282
rect 14114 29176 14148 29210
rect 14114 29104 14148 29138
rect 14114 29032 14148 29066
rect 14114 28960 14148 28994
rect 14114 28888 14148 28922
rect 14114 28816 14148 28850
rect 14114 28744 14148 28778
rect 14114 28672 14148 28706
rect 14114 28600 14148 28634
rect 14114 28528 14148 28562
rect 14114 28456 14148 28490
rect 14114 28384 14148 28418
rect 14114 28312 14148 28346
rect 14114 28240 14148 28274
rect 14114 28168 14148 28202
rect 14114 28096 14148 28130
rect 14114 28024 14148 28058
rect 14114 27952 14148 27986
rect 14114 27880 14148 27914
rect 14114 27808 14148 27842
rect 14114 27736 14148 27770
rect 14114 27664 14148 27698
rect 14114 27592 14148 27626
rect 14114 27520 14148 27554
rect 14114 27448 14148 27482
rect 14114 27376 14148 27410
rect 14114 27304 14148 27338
rect 14114 27232 14148 27266
rect 14114 27160 14148 27194
rect 14114 27088 14148 27122
rect 14114 27016 14148 27050
rect 14114 26944 14148 26978
rect 14114 26872 14148 26906
rect 14114 26800 14148 26834
rect 14114 26728 14148 26762
rect 14114 26656 14148 26690
rect 14114 26584 14148 26618
rect 14114 26512 14148 26546
rect 14114 26440 14148 26474
rect 14114 26368 14148 26402
rect 14114 26296 14148 26330
rect 14114 26224 14148 26258
rect 14114 26152 14148 26186
rect 14114 26080 14148 26114
rect 14114 26008 14148 26042
rect 14114 25936 14148 25970
rect 14114 25864 14148 25898
rect 14114 25792 14148 25826
rect 14114 25720 14148 25754
rect 14114 25648 14148 25682
rect 14114 25576 14148 25610
rect 14114 25504 14148 25538
rect 14114 25432 14148 25466
rect 14114 25360 14148 25394
rect 14114 25288 14148 25322
rect 14114 25216 14148 25250
rect 14114 25144 14148 25178
rect 14114 25072 14148 25106
rect 14114 25000 14148 25034
rect 14114 24928 14148 24962
rect 14114 24856 14148 24890
rect 14114 24784 14148 24818
rect 14114 24712 14148 24746
rect 14114 24640 14148 24674
rect 14114 24568 14148 24602
rect 14114 24496 14148 24530
rect 14114 24424 14148 24458
rect 14114 24352 14148 24386
rect 14114 24280 14148 24314
rect 14114 24208 14148 24242
rect 14114 24136 14148 24170
rect 14114 24064 14148 24098
rect 14114 23992 14148 24026
rect 14114 23920 14148 23954
rect 14114 23848 14148 23882
rect 14114 23776 14148 23810
rect 14114 23704 14148 23738
rect 14114 23632 14148 23666
rect 14114 23560 14148 23594
rect 14114 23488 14148 23522
rect 14114 23416 14148 23450
rect 14114 23344 14148 23378
rect 14114 23272 14148 23306
rect 14114 23200 14148 23234
rect 14114 23128 14148 23162
rect 14114 23056 14148 23090
rect 14114 22984 14148 23018
rect 14114 22912 14148 22946
rect 14114 22840 14148 22874
rect 14114 22768 14148 22802
rect 14114 22696 14148 22730
rect 14114 22624 14148 22658
rect 14114 22552 14148 22586
rect 14114 22480 14148 22514
rect 14114 22408 14148 22442
rect 14114 22336 14148 22370
rect 14114 22264 14148 22298
rect 14114 22192 14148 22226
rect 14114 22120 14148 22154
rect 14114 22048 14148 22082
rect 14114 21976 14148 22010
rect 14114 21904 14148 21938
rect 14114 21832 14148 21866
rect 14114 21760 14148 21794
rect 14114 21688 14148 21722
rect 14114 21616 14148 21650
rect 14114 21544 14148 21578
rect 14114 21472 14148 21506
rect 14114 21400 14148 21434
rect 14114 21328 14148 21362
rect 14114 21256 14148 21290
rect 14114 21184 14148 21218
rect 14114 21112 14148 21146
rect 14114 21040 14148 21074
rect 14114 20968 14148 21002
rect 14114 20896 14148 20930
rect 14114 20824 14148 20858
rect 14114 20752 14148 20786
rect 14114 20680 14148 20714
rect 14114 20608 14148 20642
rect 14114 20536 14148 20570
rect 14114 20464 14148 20498
rect 14114 20392 14148 20426
rect 14114 20320 14148 20354
rect 14114 20248 14148 20282
rect 14114 20176 14148 20210
rect 14114 20104 14148 20138
rect 14114 20032 14148 20066
rect 14114 19960 14148 19994
rect 14114 19888 14148 19922
rect 14114 19816 14148 19850
rect 14114 19744 14148 19778
rect 14114 19672 14148 19706
rect 14114 19600 14148 19634
rect 14114 19528 14148 19562
rect 14114 19456 14148 19490
rect 14114 19384 14148 19418
rect 14114 19312 14148 19346
rect 14114 19240 14148 19274
rect 14114 19168 14148 19202
rect 14114 19096 14148 19130
rect 14114 19024 14148 19058
rect 14114 18952 14148 18986
rect 14114 18880 14148 18914
rect 14114 18808 14148 18842
rect 14114 18736 14148 18770
rect 14114 18664 14148 18698
rect 14114 18592 14148 18626
rect 14114 18520 14148 18554
rect 14114 18448 14148 18482
rect 14114 18376 14148 18410
rect 14114 18304 14148 18338
rect 14114 18232 14148 18266
rect 14114 18160 14148 18194
rect 14114 18088 14148 18122
rect 14114 18016 14148 18050
rect 14114 17944 14148 17978
rect 14114 17872 14148 17906
rect 14114 17800 14148 17834
rect 14114 17728 14148 17762
rect 14114 17656 14148 17690
rect 14114 17584 14148 17618
rect 14114 17512 14148 17546
rect 14114 17440 14148 17474
rect 14114 17368 14148 17402
rect 14114 17296 14148 17330
rect 14114 17224 14148 17258
rect 14114 17152 14148 17186
rect 14114 17080 14148 17114
rect 14114 17008 14148 17042
rect 14114 16936 14148 16970
rect 14114 16864 14148 16898
rect 14114 16792 14148 16826
rect 14114 16720 14148 16754
rect 14114 16648 14148 16682
rect 14114 16576 14148 16610
rect 14114 16504 14148 16538
rect 14114 16432 14148 16466
rect 14114 16360 14148 16394
rect 14114 16288 14148 16322
rect 14114 16216 14148 16250
rect 14114 16144 14148 16178
rect 14114 16072 14148 16106
rect 14114 16000 14148 16034
rect 14114 15928 14148 15962
rect 14114 15856 14148 15890
rect 14114 15784 14148 15818
rect 14114 15712 14148 15746
rect 14114 15640 14148 15674
rect 14114 15568 14148 15602
rect 14114 15496 14148 15530
rect 14114 15424 14148 15458
rect 14114 15352 14148 15386
rect 14114 15280 14148 15314
rect 799 15143 833 15177
rect 799 15071 833 15105
rect 14114 15208 14148 15242
rect 14114 15136 14148 15170
rect 14114 15064 14148 15098
rect 883 14921 917 14955
rect 955 14921 989 14955
rect 1027 14921 1061 14955
rect 1099 14921 1133 14955
rect 1171 14921 1205 14955
rect 1243 14921 1277 14955
rect 1315 14921 1349 14955
rect 1387 14921 1421 14955
rect 1459 14921 1493 14955
rect 1531 14921 1565 14955
rect 1603 14921 1637 14955
rect 1675 14921 1709 14955
rect 1747 14921 1781 14955
rect 1819 14921 1853 14955
rect 1891 14921 1925 14955
rect 1963 14921 1997 14955
rect 2035 14921 2069 14955
rect 2107 14921 2141 14955
rect 2179 14921 2213 14955
rect 2251 14921 2285 14955
rect 2323 14921 2357 14955
rect 2395 14921 2429 14955
rect 2467 14921 2501 14955
rect 2539 14921 2573 14955
rect 2611 14921 2645 14955
rect 2683 14921 2717 14955
rect 2755 14921 2789 14955
rect 2827 14921 2861 14955
rect 2899 14921 2933 14955
rect 2971 14921 3005 14955
rect 3043 14921 3077 14955
rect 3115 14921 3149 14955
rect 3187 14921 3221 14955
rect 3259 14921 3293 14955
rect 3331 14921 3365 14955
rect 3403 14921 3437 14955
rect 3475 14921 3509 14955
rect 3547 14921 3581 14955
rect 3619 14921 3653 14955
rect 3691 14921 3725 14955
rect 3763 14921 3797 14955
rect 3835 14921 3869 14955
rect 3907 14921 3941 14955
rect 3979 14921 4013 14955
rect 4051 14921 4085 14955
rect 4123 14921 4157 14955
rect 4195 14921 4229 14955
rect 4267 14921 4301 14955
rect 4339 14921 4373 14955
rect 4411 14921 4445 14955
rect 4483 14921 4517 14955
rect 4555 14921 4589 14955
rect 4627 14921 4661 14955
rect 4699 14921 4733 14955
rect 4771 14921 4805 14955
rect 4843 14921 4877 14955
rect 4915 14921 4949 14955
rect 4987 14921 5021 14955
rect 5059 14921 5093 14955
rect 5131 14921 5165 14955
rect 5203 14921 5237 14955
rect 5275 14921 5309 14955
rect 5347 14921 5381 14955
rect 5419 14921 5453 14955
rect 5491 14921 5525 14955
rect 5563 14921 5597 14955
rect 5635 14921 5669 14955
rect 5707 14921 5741 14955
rect 5779 14921 5813 14955
rect 5851 14921 5885 14955
rect 5923 14921 5957 14955
rect 5995 14921 6029 14955
rect 6067 14921 6101 14955
rect 6139 14921 6173 14955
rect 6211 14921 6245 14955
rect 6283 14921 6317 14955
rect 6355 14921 6389 14955
rect 6427 14921 6461 14955
rect 6499 14921 6533 14955
rect 6571 14921 6605 14955
rect 6643 14921 6677 14955
rect 6715 14921 6749 14955
rect 6787 14921 6821 14955
rect 6859 14921 6893 14955
rect 6931 14921 6965 14955
rect 7003 14921 7037 14955
rect 7075 14921 7109 14955
rect 7147 14921 7181 14955
rect 7219 14921 7253 14955
rect 7291 14921 7325 14955
rect 7363 14921 7397 14955
rect 7435 14921 7469 14955
rect 7507 14921 7541 14955
rect 7579 14921 7613 14955
rect 7651 14921 7685 14955
rect 7723 14921 7757 14955
rect 7795 14921 7829 14955
rect 7867 14921 7901 14955
rect 7939 14921 7973 14955
rect 8011 14921 8045 14955
rect 8083 14921 8117 14955
rect 8155 14921 8189 14955
rect 8227 14921 8261 14955
rect 8299 14921 8333 14955
rect 8371 14921 8405 14955
rect 8443 14921 8477 14955
rect 8515 14921 8549 14955
rect 8587 14921 8621 14955
rect 8659 14921 8693 14955
rect 8731 14921 8765 14955
rect 8803 14921 8837 14955
rect 8875 14921 8909 14955
rect 8947 14921 8981 14955
rect 9019 14921 9053 14955
rect 9091 14921 9125 14955
rect 9163 14921 9197 14955
rect 9235 14921 9269 14955
rect 9307 14921 9341 14955
rect 9379 14921 9413 14955
rect 9451 14921 9485 14955
rect 9523 14921 9557 14955
rect 9595 14921 9629 14955
rect 9667 14921 9701 14955
rect 9739 14921 9773 14955
rect 9811 14921 9845 14955
rect 9883 14921 9917 14955
rect 9955 14921 9989 14955
rect 10027 14921 10061 14955
rect 10099 14921 10133 14955
rect 10171 14921 10205 14955
rect 10243 14921 10277 14955
rect 10315 14921 10349 14955
rect 10387 14921 10421 14955
rect 10459 14921 10493 14955
rect 10531 14921 10565 14955
rect 10603 14921 10637 14955
rect 10675 14921 10709 14955
rect 10747 14921 10781 14955
rect 10819 14921 10853 14955
rect 10891 14921 10925 14955
rect 10963 14921 10997 14955
rect 11035 14921 11069 14955
rect 11107 14921 11141 14955
rect 11179 14921 11213 14955
rect 11251 14921 11285 14955
rect 11323 14921 11357 14955
rect 11395 14921 11429 14955
rect 11467 14921 11501 14955
rect 11539 14921 11573 14955
rect 11611 14921 11645 14955
rect 11683 14921 11717 14955
rect 11755 14921 11789 14955
rect 11827 14921 11861 14955
rect 11899 14921 11933 14955
rect 11971 14921 12005 14955
rect 12043 14921 12077 14955
rect 12115 14921 12149 14955
rect 12187 14921 12221 14955
rect 12259 14921 12293 14955
rect 12331 14921 12365 14955
rect 12403 14921 12437 14955
rect 12475 14921 12509 14955
rect 12547 14921 12581 14955
rect 12619 14921 12653 14955
rect 12691 14921 12725 14955
rect 12763 14921 12797 14955
rect 12835 14921 12869 14955
rect 12907 14921 12941 14955
rect 12979 14921 13013 14955
rect 13051 14921 13085 14955
rect 13123 14921 13157 14955
rect 13195 14921 13229 14955
rect 13267 14921 13301 14955
rect 13339 14921 13373 14955
rect 13411 14921 13445 14955
rect 13483 14921 13517 14955
rect 13555 14921 13589 14955
rect 13627 14921 13661 14955
rect 13699 14921 13733 14955
rect 13771 14921 13805 14955
rect 13843 14921 13877 14955
rect 13915 14921 13949 14955
rect 13987 14921 14021 14955
rect 875 14754 894 14787
rect 894 14754 909 14787
rect 947 14754 962 14787
rect 962 14754 981 14787
rect 1019 14754 1030 14787
rect 1030 14754 1053 14787
rect 1091 14754 1098 14787
rect 1098 14754 1125 14787
rect 1163 14754 1166 14787
rect 1166 14754 1197 14787
rect 1235 14754 1268 14787
rect 1268 14754 1269 14787
rect 1307 14754 1336 14787
rect 1336 14754 1341 14787
rect 1379 14754 1404 14787
rect 1404 14754 1413 14787
rect 1451 14754 1472 14787
rect 1472 14754 1485 14787
rect 1523 14754 1540 14787
rect 1540 14754 1557 14787
rect 1595 14754 1608 14787
rect 1608 14754 1629 14787
rect 1667 14754 1676 14787
rect 1676 14754 1701 14787
rect 1739 14754 1744 14787
rect 1744 14754 1773 14787
rect 1811 14754 1812 14787
rect 1812 14754 1845 14787
rect 1883 14754 1914 14787
rect 1914 14754 1917 14787
rect 1955 14754 1982 14787
rect 1982 14754 1989 14787
rect 2027 14754 2050 14787
rect 2050 14754 2061 14787
rect 12875 14754 12896 14787
rect 12896 14754 12909 14787
rect 12947 14754 12964 14787
rect 12964 14754 12981 14787
rect 13019 14754 13032 14787
rect 13032 14754 13053 14787
rect 13091 14754 13100 14787
rect 13100 14754 13125 14787
rect 13163 14754 13168 14787
rect 13168 14754 13197 14787
rect 13235 14754 13236 14787
rect 13236 14754 13269 14787
rect 13307 14754 13338 14787
rect 13338 14754 13341 14787
rect 13379 14754 13406 14787
rect 13406 14754 13413 14787
rect 13451 14754 13474 14787
rect 13474 14754 13485 14787
rect 13523 14754 13542 14787
rect 13542 14754 13557 14787
rect 13595 14754 13610 14787
rect 13610 14754 13629 14787
rect 13667 14754 13678 14787
rect 13678 14754 13701 14787
rect 13739 14754 13746 14787
rect 13746 14754 13773 14787
rect 13811 14754 13814 14787
rect 13814 14754 13845 14787
rect 13883 14754 13916 14787
rect 13916 14754 13917 14787
rect 13955 14754 13984 14787
rect 13984 14754 13989 14787
rect 14027 14754 14052 14787
rect 14052 14754 14061 14787
rect 875 14753 909 14754
rect 947 14753 981 14754
rect 1019 14753 1053 14754
rect 1091 14753 1125 14754
rect 1163 14753 1197 14754
rect 1235 14753 1269 14754
rect 1307 14753 1341 14754
rect 1379 14753 1413 14754
rect 1451 14753 1485 14754
rect 1523 14753 1557 14754
rect 1595 14753 1629 14754
rect 1667 14753 1701 14754
rect 1739 14753 1773 14754
rect 1811 14753 1845 14754
rect 1883 14753 1917 14754
rect 1955 14753 1989 14754
rect 2027 14753 2061 14754
rect 12875 14753 12909 14754
rect 12947 14753 12981 14754
rect 13019 14753 13053 14754
rect 13091 14753 13125 14754
rect 13163 14753 13197 14754
rect 13235 14753 13269 14754
rect 13307 14753 13341 14754
rect 13379 14753 13413 14754
rect 13451 14753 13485 14754
rect 13523 14753 13557 14754
rect 13595 14753 13629 14754
rect 13667 14753 13701 14754
rect 13739 14753 13773 14754
rect 13811 14753 13845 14754
rect 13883 14753 13917 14754
rect 13955 14753 13989 14754
rect 14027 14753 14061 14754
rect 14606 36205 14633 36219
rect 14633 36205 14640 36219
rect 14606 36185 14640 36205
rect 14606 36137 14633 36147
rect 14633 36137 14640 36147
rect 14606 36113 14640 36137
rect 14606 36069 14633 36075
rect 14633 36069 14640 36075
rect 14606 36041 14640 36069
rect 14606 36001 14633 36003
rect 14633 36001 14640 36003
rect 14606 35969 14640 36001
rect 14606 35899 14640 35931
rect 14606 35897 14633 35899
rect 14633 35897 14640 35899
rect 14606 35831 14640 35859
rect 14606 35825 14633 35831
rect 14633 35825 14640 35831
rect 14606 35763 14640 35787
rect 14606 35753 14633 35763
rect 14633 35753 14640 35763
rect 14606 35695 14640 35715
rect 14606 35681 14633 35695
rect 14633 35681 14640 35695
rect 14606 35627 14640 35643
rect 14606 35609 14633 35627
rect 14633 35609 14640 35627
rect 14606 35559 14640 35571
rect 14606 35537 14633 35559
rect 14633 35537 14640 35559
rect 14606 35491 14640 35499
rect 14606 35465 14633 35491
rect 14633 35465 14640 35491
rect 14606 35423 14640 35427
rect 14606 35393 14633 35423
rect 14633 35393 14640 35423
rect 14606 35321 14633 35355
rect 14633 35321 14640 35355
rect 14606 35253 14633 35283
rect 14633 35253 14640 35283
rect 14606 35249 14640 35253
rect 14606 35185 14633 35211
rect 14633 35185 14640 35211
rect 14606 35177 14640 35185
rect 14606 35117 14633 35139
rect 14633 35117 14640 35139
rect 14606 35105 14640 35117
rect 14606 35049 14633 35067
rect 14633 35049 14640 35067
rect 14606 35033 14640 35049
rect 14606 34981 14633 34995
rect 14633 34981 14640 34995
rect 14606 34961 14640 34981
rect 14606 34913 14633 34923
rect 14633 34913 14640 34923
rect 14606 34889 14640 34913
rect 14606 34845 14633 34851
rect 14633 34845 14640 34851
rect 14606 34817 14640 34845
rect 14606 34777 14633 34779
rect 14633 34777 14640 34779
rect 14606 34745 14640 34777
rect 14606 34675 14640 34707
rect 14606 34673 14633 34675
rect 14633 34673 14640 34675
rect 14606 34607 14640 34635
rect 14606 34601 14633 34607
rect 14633 34601 14640 34607
rect 14606 34539 14640 34563
rect 14606 34529 14633 34539
rect 14633 34529 14640 34539
rect 14606 34471 14640 34491
rect 14606 34457 14633 34471
rect 14633 34457 14640 34471
rect 14606 34403 14640 34419
rect 14606 34385 14633 34403
rect 14633 34385 14640 34403
rect 14606 34335 14640 34347
rect 14606 34313 14633 34335
rect 14633 34313 14640 34335
rect 14606 34267 14640 34275
rect 14606 34241 14633 34267
rect 14633 34241 14640 34267
rect 14606 34199 14640 34203
rect 14606 34169 14633 34199
rect 14633 34169 14640 34199
rect 14606 34097 14633 34131
rect 14633 34097 14640 34131
rect 14606 34029 14633 34059
rect 14633 34029 14640 34059
rect 14606 34025 14640 34029
rect 14606 33961 14633 33987
rect 14633 33961 14640 33987
rect 14606 33953 14640 33961
rect 14606 33893 14633 33915
rect 14633 33893 14640 33915
rect 14606 33881 14640 33893
rect 14606 33825 14633 33843
rect 14633 33825 14640 33843
rect 14606 33809 14640 33825
rect 14606 33757 14633 33771
rect 14633 33757 14640 33771
rect 14606 33737 14640 33757
rect 14606 33689 14633 33699
rect 14633 33689 14640 33699
rect 14606 33665 14640 33689
rect 14606 33621 14633 33627
rect 14633 33621 14640 33627
rect 14606 33593 14640 33621
rect 14606 33553 14633 33555
rect 14633 33553 14640 33555
rect 14606 33521 14640 33553
rect 14606 33451 14640 33483
rect 14606 33449 14633 33451
rect 14633 33449 14640 33451
rect 14606 33383 14640 33411
rect 14606 33377 14633 33383
rect 14633 33377 14640 33383
rect 14606 33315 14640 33339
rect 14606 33305 14633 33315
rect 14633 33305 14640 33315
rect 14606 33247 14640 33267
rect 14606 33233 14633 33247
rect 14633 33233 14640 33247
rect 14606 33179 14640 33195
rect 14606 33161 14633 33179
rect 14633 33161 14640 33179
rect 14606 33111 14640 33123
rect 14606 33089 14633 33111
rect 14633 33089 14640 33111
rect 14606 33043 14640 33051
rect 14606 33017 14633 33043
rect 14633 33017 14640 33043
rect 14606 32975 14640 32979
rect 14606 32945 14633 32975
rect 14633 32945 14640 32975
rect 14606 32873 14633 32907
rect 14633 32873 14640 32907
rect 14606 32805 14633 32835
rect 14633 32805 14640 32835
rect 14606 32801 14640 32805
rect 14606 32737 14633 32763
rect 14633 32737 14640 32763
rect 14606 32729 14640 32737
rect 14606 32669 14633 32691
rect 14633 32669 14640 32691
rect 14606 32657 14640 32669
rect 14606 32601 14633 32619
rect 14633 32601 14640 32619
rect 14606 32585 14640 32601
rect 14606 32533 14633 32547
rect 14633 32533 14640 32547
rect 14606 32513 14640 32533
rect 14606 32465 14633 32475
rect 14633 32465 14640 32475
rect 14606 32441 14640 32465
rect 14606 32397 14633 32403
rect 14633 32397 14640 32403
rect 14606 32369 14640 32397
rect 14606 32329 14633 32331
rect 14633 32329 14640 32331
rect 14606 32297 14640 32329
rect 14606 32227 14640 32259
rect 14606 32225 14633 32227
rect 14633 32225 14640 32227
rect 14606 32159 14640 32187
rect 14606 32153 14633 32159
rect 14633 32153 14640 32159
rect 14606 32091 14640 32115
rect 14606 32081 14633 32091
rect 14633 32081 14640 32091
rect 14606 32023 14640 32043
rect 14606 32009 14633 32023
rect 14633 32009 14640 32023
rect 14606 31955 14640 31971
rect 14606 31937 14633 31955
rect 14633 31937 14640 31955
rect 14606 31887 14640 31899
rect 14606 31865 14633 31887
rect 14633 31865 14640 31887
rect 14606 31819 14640 31827
rect 14606 31793 14633 31819
rect 14633 31793 14640 31819
rect 14606 31751 14640 31755
rect 14606 31721 14633 31751
rect 14633 31721 14640 31751
rect 14606 31649 14633 31683
rect 14633 31649 14640 31683
rect 14606 31581 14633 31611
rect 14633 31581 14640 31611
rect 14606 31577 14640 31581
rect 14606 31513 14633 31539
rect 14633 31513 14640 31539
rect 14606 31505 14640 31513
rect 14606 31445 14633 31467
rect 14633 31445 14640 31467
rect 14606 31433 14640 31445
rect 14606 31377 14633 31395
rect 14633 31377 14640 31395
rect 14606 31361 14640 31377
rect 14606 31309 14633 31323
rect 14633 31309 14640 31323
rect 14606 31289 14640 31309
rect 14606 31241 14633 31251
rect 14633 31241 14640 31251
rect 14606 31217 14640 31241
rect 14606 31173 14633 31179
rect 14633 31173 14640 31179
rect 14606 31145 14640 31173
rect 14606 31105 14633 31107
rect 14633 31105 14640 31107
rect 14606 31073 14640 31105
rect 14606 31003 14640 31035
rect 14606 31001 14633 31003
rect 14633 31001 14640 31003
rect 14606 30935 14640 30963
rect 14606 30929 14633 30935
rect 14633 30929 14640 30935
rect 14606 30867 14640 30891
rect 14606 30857 14633 30867
rect 14633 30857 14640 30867
rect 14606 30799 14640 30819
rect 14606 30785 14633 30799
rect 14633 30785 14640 30799
rect 14606 30731 14640 30747
rect 14606 30713 14633 30731
rect 14633 30713 14640 30731
rect 14606 30663 14640 30675
rect 14606 30641 14633 30663
rect 14633 30641 14640 30663
rect 14606 30595 14640 30603
rect 14606 30569 14633 30595
rect 14633 30569 14640 30595
rect 14606 30527 14640 30531
rect 14606 30497 14633 30527
rect 14633 30497 14640 30527
rect 14606 30425 14633 30459
rect 14633 30425 14640 30459
rect 14606 30357 14633 30387
rect 14633 30357 14640 30387
rect 14606 30353 14640 30357
rect 14606 30289 14633 30315
rect 14633 30289 14640 30315
rect 14606 30281 14640 30289
rect 14606 30221 14633 30243
rect 14633 30221 14640 30243
rect 14606 30209 14640 30221
rect 14606 30153 14633 30171
rect 14633 30153 14640 30171
rect 14606 30137 14640 30153
rect 14606 30085 14633 30099
rect 14633 30085 14640 30099
rect 14606 30065 14640 30085
rect 14606 30017 14633 30027
rect 14633 30017 14640 30027
rect 14606 29993 14640 30017
rect 14606 29949 14633 29955
rect 14633 29949 14640 29955
rect 14606 29921 14640 29949
rect 14606 29881 14633 29883
rect 14633 29881 14640 29883
rect 14606 29849 14640 29881
rect 14606 29779 14640 29811
rect 14606 29777 14633 29779
rect 14633 29777 14640 29779
rect 14606 29711 14640 29739
rect 14606 29705 14633 29711
rect 14633 29705 14640 29711
rect 14606 29643 14640 29667
rect 14606 29633 14633 29643
rect 14633 29633 14640 29643
rect 14606 29575 14640 29595
rect 14606 29561 14633 29575
rect 14633 29561 14640 29575
rect 14606 29507 14640 29523
rect 14606 29489 14633 29507
rect 14633 29489 14640 29507
rect 14606 29439 14640 29451
rect 14606 29417 14633 29439
rect 14633 29417 14640 29439
rect 14606 29371 14640 29379
rect 14606 29345 14633 29371
rect 14633 29345 14640 29371
rect 14606 29303 14640 29307
rect 14606 29273 14633 29303
rect 14633 29273 14640 29303
rect 14606 29201 14633 29235
rect 14633 29201 14640 29235
rect 14606 29133 14633 29163
rect 14633 29133 14640 29163
rect 14606 29129 14640 29133
rect 14606 29065 14633 29091
rect 14633 29065 14640 29091
rect 14606 29057 14640 29065
rect 14606 28997 14633 29019
rect 14633 28997 14640 29019
rect 14606 28985 14640 28997
rect 14606 28929 14633 28947
rect 14633 28929 14640 28947
rect 14606 28913 14640 28929
rect 14606 28861 14633 28875
rect 14633 28861 14640 28875
rect 14606 28841 14640 28861
rect 14606 28793 14633 28803
rect 14633 28793 14640 28803
rect 14606 28769 14640 28793
rect 14606 28725 14633 28731
rect 14633 28725 14640 28731
rect 14606 28697 14640 28725
rect 14606 28657 14633 28659
rect 14633 28657 14640 28659
rect 14606 28625 14640 28657
rect 14606 28555 14640 28587
rect 14606 28553 14633 28555
rect 14633 28553 14640 28555
rect 14606 28487 14640 28515
rect 14606 28481 14633 28487
rect 14633 28481 14640 28487
rect 14606 28419 14640 28443
rect 14606 28409 14633 28419
rect 14633 28409 14640 28419
rect 14606 28351 14640 28371
rect 14606 28337 14633 28351
rect 14633 28337 14640 28351
rect 14606 28283 14640 28299
rect 14606 28265 14633 28283
rect 14633 28265 14640 28283
rect 14606 28215 14640 28227
rect 14606 28193 14633 28215
rect 14633 28193 14640 28215
rect 14606 28147 14640 28155
rect 14606 28121 14633 28147
rect 14633 28121 14640 28147
rect 14606 28079 14640 28083
rect 14606 28049 14633 28079
rect 14633 28049 14640 28079
rect 14606 27977 14633 28011
rect 14633 27977 14640 28011
rect 14606 27909 14633 27939
rect 14633 27909 14640 27939
rect 14606 27905 14640 27909
rect 14606 27841 14633 27867
rect 14633 27841 14640 27867
rect 14606 27833 14640 27841
rect 14606 27773 14633 27795
rect 14633 27773 14640 27795
rect 14606 27761 14640 27773
rect 14606 27705 14633 27723
rect 14633 27705 14640 27723
rect 14606 27689 14640 27705
rect 14606 27637 14633 27651
rect 14633 27637 14640 27651
rect 14606 27617 14640 27637
rect 14606 27569 14633 27579
rect 14633 27569 14640 27579
rect 14606 27545 14640 27569
rect 14606 27501 14633 27507
rect 14633 27501 14640 27507
rect 14606 27473 14640 27501
rect 14606 27433 14633 27435
rect 14633 27433 14640 27435
rect 14606 27401 14640 27433
rect 14606 27331 14640 27363
rect 14606 27329 14633 27331
rect 14633 27329 14640 27331
rect 14606 27263 14640 27291
rect 14606 27257 14633 27263
rect 14633 27257 14640 27263
rect 14606 27195 14640 27219
rect 14606 27185 14633 27195
rect 14633 27185 14640 27195
rect 14606 27127 14640 27147
rect 14606 27113 14633 27127
rect 14633 27113 14640 27127
rect 14606 27059 14640 27075
rect 14606 27041 14633 27059
rect 14633 27041 14640 27059
rect 14606 26991 14640 27003
rect 14606 26969 14633 26991
rect 14633 26969 14640 26991
rect 14606 26923 14640 26931
rect 14606 26897 14633 26923
rect 14633 26897 14640 26923
rect 14606 26855 14640 26859
rect 14606 26825 14633 26855
rect 14633 26825 14640 26855
rect 14606 26753 14633 26787
rect 14633 26753 14640 26787
rect 14606 26685 14633 26715
rect 14633 26685 14640 26715
rect 14606 26681 14640 26685
rect 14606 26617 14633 26643
rect 14633 26617 14640 26643
rect 14606 26609 14640 26617
rect 14606 26549 14633 26571
rect 14633 26549 14640 26571
rect 14606 26537 14640 26549
rect 14606 26481 14633 26499
rect 14633 26481 14640 26499
rect 14606 26465 14640 26481
rect 14606 26413 14633 26427
rect 14633 26413 14640 26427
rect 14606 26393 14640 26413
rect 14606 26345 14633 26355
rect 14633 26345 14640 26355
rect 14606 26321 14640 26345
rect 14606 26277 14633 26283
rect 14633 26277 14640 26283
rect 14606 26249 14640 26277
rect 14606 26209 14633 26211
rect 14633 26209 14640 26211
rect 14606 26177 14640 26209
rect 14606 26107 14640 26139
rect 14606 26105 14633 26107
rect 14633 26105 14640 26107
rect 14606 26039 14640 26067
rect 14606 26033 14633 26039
rect 14633 26033 14640 26039
rect 14606 25971 14640 25995
rect 14606 25961 14633 25971
rect 14633 25961 14640 25971
rect 14606 25903 14640 25923
rect 14606 25889 14633 25903
rect 14633 25889 14640 25903
rect 14606 25835 14640 25851
rect 14606 25817 14633 25835
rect 14633 25817 14640 25835
rect 14606 25767 14640 25779
rect 14606 25745 14633 25767
rect 14633 25745 14640 25767
rect 14606 25699 14640 25707
rect 14606 25673 14633 25699
rect 14633 25673 14640 25699
rect 14606 25631 14640 25635
rect 14606 25601 14633 25631
rect 14633 25601 14640 25631
rect 14606 25529 14633 25563
rect 14633 25529 14640 25563
rect 14606 25461 14633 25491
rect 14633 25461 14640 25491
rect 14606 25457 14640 25461
rect 14606 25393 14633 25419
rect 14633 25393 14640 25419
rect 14606 25385 14640 25393
rect 14606 25325 14633 25347
rect 14633 25325 14640 25347
rect 14606 25313 14640 25325
rect 14606 25257 14633 25275
rect 14633 25257 14640 25275
rect 14606 25241 14640 25257
rect 14606 25189 14633 25203
rect 14633 25189 14640 25203
rect 14606 25169 14640 25189
rect 14606 25121 14633 25131
rect 14633 25121 14640 25131
rect 14606 25097 14640 25121
rect 14606 25053 14633 25059
rect 14633 25053 14640 25059
rect 14606 25025 14640 25053
rect 14606 24985 14633 24987
rect 14633 24985 14640 24987
rect 14606 24953 14640 24985
rect 14606 24883 14640 24915
rect 14606 24881 14633 24883
rect 14633 24881 14640 24883
rect 14606 24815 14640 24843
rect 14606 24809 14633 24815
rect 14633 24809 14640 24815
rect 14606 24747 14640 24771
rect 14606 24737 14633 24747
rect 14633 24737 14640 24747
rect 14606 24679 14640 24699
rect 14606 24665 14633 24679
rect 14633 24665 14640 24679
rect 14606 24611 14640 24627
rect 14606 24593 14633 24611
rect 14633 24593 14640 24611
rect 14606 24543 14640 24555
rect 14606 24521 14633 24543
rect 14633 24521 14640 24543
rect 14606 24475 14640 24483
rect 14606 24449 14633 24475
rect 14633 24449 14640 24475
rect 14606 24407 14640 24411
rect 14606 24377 14633 24407
rect 14633 24377 14640 24407
rect 14606 24305 14633 24339
rect 14633 24305 14640 24339
rect 14606 24237 14633 24267
rect 14633 24237 14640 24267
rect 14606 24233 14640 24237
rect 14606 24169 14633 24195
rect 14633 24169 14640 24195
rect 14606 24161 14640 24169
rect 14606 24101 14633 24123
rect 14633 24101 14640 24123
rect 14606 24089 14640 24101
rect 14606 24033 14633 24051
rect 14633 24033 14640 24051
rect 14606 24017 14640 24033
rect 14606 23965 14633 23979
rect 14633 23965 14640 23979
rect 14606 23945 14640 23965
rect 14606 23897 14633 23907
rect 14633 23897 14640 23907
rect 14606 23873 14640 23897
rect 14606 23829 14633 23835
rect 14633 23829 14640 23835
rect 14606 23801 14640 23829
rect 14606 23761 14633 23763
rect 14633 23761 14640 23763
rect 14606 23729 14640 23761
rect 14606 23659 14640 23691
rect 14606 23657 14633 23659
rect 14633 23657 14640 23659
rect 14606 23591 14640 23619
rect 14606 23585 14633 23591
rect 14633 23585 14640 23591
rect 14606 23523 14640 23547
rect 14606 23513 14633 23523
rect 14633 23513 14640 23523
rect 14606 23455 14640 23475
rect 14606 23441 14633 23455
rect 14633 23441 14640 23455
rect 14606 23387 14640 23403
rect 14606 23369 14633 23387
rect 14633 23369 14640 23387
rect 14606 23319 14640 23331
rect 14606 23297 14633 23319
rect 14633 23297 14640 23319
rect 14606 23251 14640 23259
rect 14606 23225 14633 23251
rect 14633 23225 14640 23251
rect 14606 23183 14640 23187
rect 14606 23153 14633 23183
rect 14633 23153 14640 23183
rect 14606 23081 14633 23115
rect 14633 23081 14640 23115
rect 14606 23013 14633 23043
rect 14633 23013 14640 23043
rect 14606 23009 14640 23013
rect 14606 22945 14633 22971
rect 14633 22945 14640 22971
rect 14606 22937 14640 22945
rect 14606 22877 14633 22899
rect 14633 22877 14640 22899
rect 14606 22865 14640 22877
rect 14606 22809 14633 22827
rect 14633 22809 14640 22827
rect 14606 22793 14640 22809
rect 14606 22741 14633 22755
rect 14633 22741 14640 22755
rect 14606 22721 14640 22741
rect 14606 22673 14633 22683
rect 14633 22673 14640 22683
rect 14606 22649 14640 22673
rect 14606 22605 14633 22611
rect 14633 22605 14640 22611
rect 14606 22577 14640 22605
rect 14606 22537 14633 22539
rect 14633 22537 14640 22539
rect 14606 22505 14640 22537
rect 14606 22435 14640 22467
rect 14606 22433 14633 22435
rect 14633 22433 14640 22435
rect 14606 22367 14640 22395
rect 14606 22361 14633 22367
rect 14633 22361 14640 22367
rect 14606 22299 14640 22323
rect 14606 22289 14633 22299
rect 14633 22289 14640 22299
rect 14606 22231 14640 22251
rect 14606 22217 14633 22231
rect 14633 22217 14640 22231
rect 14606 22163 14640 22179
rect 14606 22145 14633 22163
rect 14633 22145 14640 22163
rect 14606 22095 14640 22107
rect 14606 22073 14633 22095
rect 14633 22073 14640 22095
rect 14606 22027 14640 22035
rect 14606 22001 14633 22027
rect 14633 22001 14640 22027
rect 14606 21959 14640 21963
rect 14606 21929 14633 21959
rect 14633 21929 14640 21959
rect 14606 21857 14633 21891
rect 14633 21857 14640 21891
rect 14606 21789 14633 21819
rect 14633 21789 14640 21819
rect 14606 21785 14640 21789
rect 14606 21721 14633 21747
rect 14633 21721 14640 21747
rect 14606 21713 14640 21721
rect 14606 21653 14633 21675
rect 14633 21653 14640 21675
rect 14606 21641 14640 21653
rect 14606 21585 14633 21603
rect 14633 21585 14640 21603
rect 14606 21569 14640 21585
rect 14606 21517 14633 21531
rect 14633 21517 14640 21531
rect 14606 21497 14640 21517
rect 14606 21449 14633 21459
rect 14633 21449 14640 21459
rect 14606 21425 14640 21449
rect 14606 21381 14633 21387
rect 14633 21381 14640 21387
rect 14606 21353 14640 21381
rect 14606 21313 14633 21315
rect 14633 21313 14640 21315
rect 14606 21281 14640 21313
rect 14606 21211 14640 21243
rect 14606 21209 14633 21211
rect 14633 21209 14640 21211
rect 14606 21143 14640 21171
rect 14606 21137 14633 21143
rect 14633 21137 14640 21143
rect 14606 21075 14640 21099
rect 14606 21065 14633 21075
rect 14633 21065 14640 21075
rect 14606 21007 14640 21027
rect 14606 20993 14633 21007
rect 14633 20993 14640 21007
rect 14606 20939 14640 20955
rect 14606 20921 14633 20939
rect 14633 20921 14640 20939
rect 14606 20871 14640 20883
rect 14606 20849 14633 20871
rect 14633 20849 14640 20871
rect 14606 20803 14640 20811
rect 14606 20777 14633 20803
rect 14633 20777 14640 20803
rect 14606 20735 14640 20739
rect 14606 20705 14633 20735
rect 14633 20705 14640 20735
rect 14606 20633 14633 20667
rect 14633 20633 14640 20667
rect 14606 20565 14633 20595
rect 14633 20565 14640 20595
rect 14606 20561 14640 20565
rect 14606 20497 14633 20523
rect 14633 20497 14640 20523
rect 14606 20489 14640 20497
rect 14606 20429 14633 20451
rect 14633 20429 14640 20451
rect 14606 20417 14640 20429
rect 14606 20361 14633 20379
rect 14633 20361 14640 20379
rect 14606 20345 14640 20361
rect 14606 20293 14633 20307
rect 14633 20293 14640 20307
rect 14606 20273 14640 20293
rect 14606 20225 14633 20235
rect 14633 20225 14640 20235
rect 14606 20201 14640 20225
rect 14606 20157 14633 20163
rect 14633 20157 14640 20163
rect 14606 20129 14640 20157
rect 14606 20089 14633 20091
rect 14633 20089 14640 20091
rect 14606 20057 14640 20089
rect 14606 19987 14640 20019
rect 14606 19985 14633 19987
rect 14633 19985 14640 19987
rect 14606 19919 14640 19947
rect 14606 19913 14633 19919
rect 14633 19913 14640 19919
rect 14606 19851 14640 19875
rect 14606 19841 14633 19851
rect 14633 19841 14640 19851
rect 14606 19783 14640 19803
rect 14606 19769 14633 19783
rect 14633 19769 14640 19783
rect 14606 19715 14640 19731
rect 14606 19697 14633 19715
rect 14633 19697 14640 19715
rect 14606 19647 14640 19659
rect 14606 19625 14633 19647
rect 14633 19625 14640 19647
rect 14606 19579 14640 19587
rect 14606 19553 14633 19579
rect 14633 19553 14640 19579
rect 14606 19511 14640 19515
rect 14606 19481 14633 19511
rect 14633 19481 14640 19511
rect 14606 19409 14633 19443
rect 14633 19409 14640 19443
rect 14606 19341 14633 19371
rect 14633 19341 14640 19371
rect 14606 19337 14640 19341
rect 14606 19273 14633 19299
rect 14633 19273 14640 19299
rect 14606 19265 14640 19273
rect 14606 19205 14633 19227
rect 14633 19205 14640 19227
rect 14606 19193 14640 19205
rect 14606 19137 14633 19155
rect 14633 19137 14640 19155
rect 14606 19121 14640 19137
rect 14606 19069 14633 19083
rect 14633 19069 14640 19083
rect 14606 19049 14640 19069
rect 14606 19001 14633 19011
rect 14633 19001 14640 19011
rect 14606 18977 14640 19001
rect 14606 18933 14633 18939
rect 14633 18933 14640 18939
rect 14606 18905 14640 18933
rect 14606 18865 14633 18867
rect 14633 18865 14640 18867
rect 14606 18833 14640 18865
rect 14606 18763 14640 18795
rect 14606 18761 14633 18763
rect 14633 18761 14640 18763
rect 14606 18695 14640 18723
rect 14606 18689 14633 18695
rect 14633 18689 14640 18695
rect 14606 18627 14640 18651
rect 14606 18617 14633 18627
rect 14633 18617 14640 18627
rect 14606 18559 14640 18579
rect 14606 18545 14633 18559
rect 14633 18545 14640 18559
rect 14606 18491 14640 18507
rect 14606 18473 14633 18491
rect 14633 18473 14640 18491
rect 14606 18423 14640 18435
rect 14606 18401 14633 18423
rect 14633 18401 14640 18423
rect 14606 18355 14640 18363
rect 14606 18329 14633 18355
rect 14633 18329 14640 18355
rect 14606 18287 14640 18291
rect 14606 18257 14633 18287
rect 14633 18257 14640 18287
rect 14606 18185 14633 18219
rect 14633 18185 14640 18219
rect 14606 18117 14633 18147
rect 14633 18117 14640 18147
rect 14606 18113 14640 18117
rect 14606 18049 14633 18075
rect 14633 18049 14640 18075
rect 14606 18041 14640 18049
rect 14606 17981 14633 18003
rect 14633 17981 14640 18003
rect 14606 17969 14640 17981
rect 14606 17913 14633 17931
rect 14633 17913 14640 17931
rect 14606 17897 14640 17913
rect 14606 17845 14633 17859
rect 14633 17845 14640 17859
rect 14606 17825 14640 17845
rect 14606 17777 14633 17787
rect 14633 17777 14640 17787
rect 14606 17753 14640 17777
rect 14606 17709 14633 17715
rect 14633 17709 14640 17715
rect 14606 17681 14640 17709
rect 14606 17641 14633 17643
rect 14633 17641 14640 17643
rect 14606 17609 14640 17641
rect 14606 17539 14640 17571
rect 14606 17537 14633 17539
rect 14633 17537 14640 17539
rect 14606 17471 14640 17499
rect 14606 17465 14633 17471
rect 14633 17465 14640 17471
rect 14606 17403 14640 17427
rect 14606 17393 14633 17403
rect 14633 17393 14640 17403
rect 14606 17335 14640 17355
rect 14606 17321 14633 17335
rect 14633 17321 14640 17335
rect 14606 17267 14640 17283
rect 14606 17249 14633 17267
rect 14633 17249 14640 17267
rect 14606 17199 14640 17211
rect 14606 17177 14633 17199
rect 14633 17177 14640 17199
rect 14606 17131 14640 17139
rect 14606 17105 14633 17131
rect 14633 17105 14640 17131
rect 14606 17063 14640 17067
rect 14606 17033 14633 17063
rect 14633 17033 14640 17063
rect 14606 16961 14633 16995
rect 14633 16961 14640 16995
rect 14606 16893 14633 16923
rect 14633 16893 14640 16923
rect 14606 16889 14640 16893
rect 14606 16825 14633 16851
rect 14633 16825 14640 16851
rect 14606 16817 14640 16825
rect 14606 16757 14633 16779
rect 14633 16757 14640 16779
rect 14606 16745 14640 16757
rect 14606 16689 14633 16707
rect 14633 16689 14640 16707
rect 14606 16673 14640 16689
rect 14606 16621 14633 16635
rect 14633 16621 14640 16635
rect 14606 16601 14640 16621
rect 14606 16553 14633 16563
rect 14633 16553 14640 16563
rect 14606 16529 14640 16553
rect 14606 16485 14633 16491
rect 14633 16485 14640 16491
rect 14606 16457 14640 16485
rect 14606 16417 14633 16419
rect 14633 16417 14640 16419
rect 14606 16385 14640 16417
rect 14606 16315 14640 16347
rect 14606 16313 14633 16315
rect 14633 16313 14640 16315
rect 14606 16247 14640 16275
rect 14606 16241 14633 16247
rect 14633 16241 14640 16247
rect 14606 16179 14640 16203
rect 14606 16169 14633 16179
rect 14633 16169 14640 16179
rect 14606 16111 14640 16131
rect 14606 16097 14633 16111
rect 14633 16097 14640 16111
rect 14606 16043 14640 16059
rect 14606 16025 14633 16043
rect 14633 16025 14640 16043
rect 14606 15975 14640 15987
rect 14606 15953 14633 15975
rect 14633 15953 14640 15975
rect 14606 15907 14640 15915
rect 14606 15881 14633 15907
rect 14633 15881 14640 15907
rect 14606 15839 14640 15843
rect 14606 15809 14633 15839
rect 14633 15809 14640 15839
rect 14606 15737 14633 15771
rect 14633 15737 14640 15771
rect 14606 15669 14633 15699
rect 14633 15669 14640 15699
rect 14606 15665 14640 15669
rect 14606 15601 14633 15627
rect 14633 15601 14640 15627
rect 14606 15593 14640 15601
rect 14606 15533 14633 15555
rect 14633 15533 14640 15555
rect 14606 15521 14640 15533
rect 14606 15465 14633 15483
rect 14633 15465 14640 15483
rect 14606 15449 14640 15465
rect 14606 15397 14633 15411
rect 14633 15397 14640 15411
rect 14606 15377 14640 15397
rect 14606 15329 14633 15339
rect 14633 15329 14640 15339
rect 14606 15305 14640 15329
rect 14606 15261 14633 15267
rect 14633 15261 14640 15267
rect 14606 15233 14640 15261
rect 14606 15193 14633 15195
rect 14633 15193 14640 15195
rect 14606 15161 14640 15193
rect 14606 15091 14640 15123
rect 14606 15089 14633 15091
rect 14633 15089 14640 15091
rect 14606 15023 14640 15051
rect 14606 15017 14633 15023
rect 14633 15017 14640 15023
rect 14606 14955 14640 14979
rect 14606 14945 14633 14955
rect 14633 14945 14640 14955
rect 14606 14887 14640 14907
rect 14606 14873 14633 14887
rect 14633 14873 14640 14887
rect 14606 14819 14640 14835
rect 14606 14801 14633 14819
rect 14633 14801 14640 14819
rect 14606 14751 14640 14763
rect 312 14677 346 14694
rect 312 14660 338 14677
rect 338 14660 346 14677
rect 14606 14729 14633 14751
rect 14633 14729 14640 14751
rect 14606 14683 14640 14691
rect 14606 14657 14633 14683
rect 14633 14657 14640 14683
rect 312 14431 346 14465
rect 602 14464 636 14465
rect 2303 14464 2337 14465
rect 2375 14464 2409 14465
rect 2447 14464 2481 14465
rect 2519 14464 2553 14465
rect 2591 14464 2625 14465
rect 2663 14464 2697 14465
rect 2735 14464 2769 14465
rect 2807 14464 2841 14465
rect 2879 14464 2913 14465
rect 2951 14464 2985 14465
rect 3023 14464 3057 14465
rect 3095 14464 3129 14465
rect 3167 14464 3201 14465
rect 3239 14464 3273 14465
rect 3311 14464 3345 14465
rect 3383 14464 3417 14465
rect 3455 14464 3489 14465
rect 3527 14464 3561 14465
rect 3599 14464 3633 14465
rect 3671 14464 3705 14465
rect 3743 14464 3777 14465
rect 3815 14464 3849 14465
rect 3887 14464 3921 14465
rect 3959 14464 3993 14465
rect 4031 14464 4065 14465
rect 4103 14464 4137 14465
rect 4175 14464 4209 14465
rect 4247 14464 4281 14465
rect 4319 14464 4353 14465
rect 4391 14464 4425 14465
rect 4463 14464 4497 14465
rect 4535 14464 4569 14465
rect 4607 14464 4641 14465
rect 4679 14464 4713 14465
rect 4751 14464 4785 14465
rect 4823 14464 4857 14465
rect 4895 14464 4929 14465
rect 4967 14464 5001 14465
rect 5039 14464 5073 14465
rect 5111 14464 5145 14465
rect 5183 14464 5217 14465
rect 5255 14464 5289 14465
rect 5327 14464 5361 14465
rect 5399 14464 5433 14465
rect 5471 14464 5505 14465
rect 5543 14464 5577 14465
rect 5615 14464 5649 14465
rect 5687 14464 5721 14465
rect 5759 14464 5793 14465
rect 5831 14464 5865 14465
rect 5903 14464 5937 14465
rect 5975 14464 6009 14465
rect 6047 14464 6081 14465
rect 6119 14464 6153 14465
rect 6191 14464 6225 14465
rect 6263 14464 6297 14465
rect 6335 14464 6369 14465
rect 6407 14464 6441 14465
rect 6479 14464 6513 14465
rect 6551 14464 6585 14465
rect 6623 14464 6657 14465
rect 6695 14464 6729 14465
rect 6767 14464 6801 14465
rect 6839 14464 6873 14465
rect 6911 14464 6945 14465
rect 6983 14464 7017 14465
rect 7055 14464 7089 14465
rect 7127 14464 7161 14465
rect 7199 14464 7233 14465
rect 7271 14464 7305 14465
rect 7343 14464 7377 14465
rect 7415 14464 7449 14465
rect 7487 14464 7521 14465
rect 7559 14464 7593 14465
rect 7631 14464 7665 14465
rect 7703 14464 7737 14465
rect 7775 14464 7809 14465
rect 7847 14464 7881 14465
rect 7919 14464 7953 14465
rect 7991 14464 8025 14465
rect 8063 14464 8097 14465
rect 8135 14464 8169 14465
rect 8207 14464 8241 14465
rect 8279 14464 8313 14465
rect 8351 14464 8385 14465
rect 8423 14464 8457 14465
rect 8495 14464 8529 14465
rect 8567 14464 8601 14465
rect 8639 14464 8673 14465
rect 8711 14464 8745 14465
rect 8783 14464 8817 14465
rect 8855 14464 8889 14465
rect 8927 14464 8961 14465
rect 8999 14464 9033 14465
rect 9071 14464 9105 14465
rect 9143 14464 9177 14465
rect 9215 14464 9249 14465
rect 9287 14464 9321 14465
rect 9359 14464 9393 14465
rect 9431 14464 9465 14465
rect 9503 14464 9537 14465
rect 9575 14464 9609 14465
rect 9647 14464 9681 14465
rect 9719 14464 9753 14465
rect 9791 14464 9825 14465
rect 9863 14464 9897 14465
rect 9935 14464 9969 14465
rect 10007 14464 10041 14465
rect 10079 14464 10113 14465
rect 10151 14464 10185 14465
rect 10223 14464 10257 14465
rect 10295 14464 10329 14465
rect 10367 14464 10401 14465
rect 10439 14464 10473 14465
rect 10511 14464 10545 14465
rect 10583 14464 10617 14465
rect 10655 14464 10689 14465
rect 10727 14464 10761 14465
rect 10799 14464 10833 14465
rect 10871 14464 10905 14465
rect 10943 14464 10977 14465
rect 11015 14464 11049 14465
rect 11087 14464 11121 14465
rect 11159 14464 11193 14465
rect 11231 14464 11265 14465
rect 11303 14464 11337 14465
rect 11375 14464 11409 14465
rect 11447 14464 11481 14465
rect 11519 14464 11553 14465
rect 11591 14464 11625 14465
rect 11663 14464 11697 14465
rect 11735 14464 11769 14465
rect 11807 14464 11841 14465
rect 11879 14464 11913 14465
rect 11951 14464 11985 14465
rect 12023 14464 12057 14465
rect 12095 14464 12129 14465
rect 12167 14464 12201 14465
rect 12239 14464 12273 14465
rect 12311 14464 12345 14465
rect 12383 14464 12417 14465
rect 12455 14464 12489 14465
rect 12527 14464 12561 14465
rect 12599 14464 12633 14465
rect 602 14431 604 14464
rect 604 14431 636 14464
rect 2303 14431 2304 14464
rect 2304 14431 2337 14464
rect 2375 14431 2406 14464
rect 2406 14431 2409 14464
rect 2447 14431 2474 14464
rect 2474 14431 2481 14464
rect 2519 14431 2542 14464
rect 2542 14431 2553 14464
rect 2591 14431 2610 14464
rect 2610 14431 2625 14464
rect 2663 14431 2678 14464
rect 2678 14431 2697 14464
rect 2735 14431 2746 14464
rect 2746 14431 2769 14464
rect 2807 14431 2814 14464
rect 2814 14431 2841 14464
rect 2879 14431 2882 14464
rect 2882 14431 2913 14464
rect 2951 14431 2984 14464
rect 2984 14431 2985 14464
rect 3023 14431 3052 14464
rect 3052 14431 3057 14464
rect 3095 14431 3120 14464
rect 3120 14431 3129 14464
rect 3167 14431 3188 14464
rect 3188 14431 3201 14464
rect 3239 14431 3256 14464
rect 3256 14431 3273 14464
rect 3311 14431 3324 14464
rect 3324 14431 3345 14464
rect 3383 14431 3392 14464
rect 3392 14431 3417 14464
rect 3455 14431 3460 14464
rect 3460 14431 3489 14464
rect 3527 14431 3528 14464
rect 3528 14431 3561 14464
rect 3599 14431 3630 14464
rect 3630 14431 3633 14464
rect 3671 14431 3698 14464
rect 3698 14431 3705 14464
rect 3743 14431 3766 14464
rect 3766 14431 3777 14464
rect 3815 14431 3834 14464
rect 3834 14431 3849 14464
rect 3887 14431 3902 14464
rect 3902 14431 3921 14464
rect 3959 14431 3970 14464
rect 3970 14431 3993 14464
rect 4031 14431 4038 14464
rect 4038 14431 4065 14464
rect 4103 14431 4106 14464
rect 4106 14431 4137 14464
rect 4175 14431 4208 14464
rect 4208 14431 4209 14464
rect 4247 14431 4276 14464
rect 4276 14431 4281 14464
rect 4319 14431 4344 14464
rect 4344 14431 4353 14464
rect 4391 14431 4412 14464
rect 4412 14431 4425 14464
rect 4463 14431 4480 14464
rect 4480 14431 4497 14464
rect 4535 14431 4548 14464
rect 4548 14431 4569 14464
rect 4607 14431 4616 14464
rect 4616 14431 4641 14464
rect 4679 14431 4684 14464
rect 4684 14431 4713 14464
rect 4751 14431 4752 14464
rect 4752 14431 4785 14464
rect 4823 14431 4854 14464
rect 4854 14431 4857 14464
rect 4895 14431 4922 14464
rect 4922 14431 4929 14464
rect 4967 14431 4990 14464
rect 4990 14431 5001 14464
rect 5039 14431 5058 14464
rect 5058 14431 5073 14464
rect 5111 14431 5126 14464
rect 5126 14431 5145 14464
rect 5183 14431 5194 14464
rect 5194 14431 5217 14464
rect 5255 14431 5262 14464
rect 5262 14431 5289 14464
rect 5327 14431 5330 14464
rect 5330 14431 5361 14464
rect 5399 14431 5432 14464
rect 5432 14431 5433 14464
rect 5471 14431 5500 14464
rect 5500 14431 5505 14464
rect 5543 14431 5568 14464
rect 5568 14431 5577 14464
rect 5615 14431 5636 14464
rect 5636 14431 5649 14464
rect 5687 14431 5704 14464
rect 5704 14431 5721 14464
rect 5759 14431 5772 14464
rect 5772 14431 5793 14464
rect 5831 14431 5840 14464
rect 5840 14431 5865 14464
rect 5903 14431 5908 14464
rect 5908 14431 5937 14464
rect 5975 14431 5976 14464
rect 5976 14431 6009 14464
rect 6047 14431 6078 14464
rect 6078 14431 6081 14464
rect 6119 14431 6146 14464
rect 6146 14431 6153 14464
rect 6191 14431 6214 14464
rect 6214 14431 6225 14464
rect 6263 14431 6282 14464
rect 6282 14431 6297 14464
rect 6335 14431 6350 14464
rect 6350 14431 6369 14464
rect 6407 14431 6418 14464
rect 6418 14431 6441 14464
rect 6479 14431 6486 14464
rect 6486 14431 6513 14464
rect 6551 14431 6554 14464
rect 6554 14431 6585 14464
rect 6623 14431 6656 14464
rect 6656 14431 6657 14464
rect 6695 14431 6724 14464
rect 6724 14431 6729 14464
rect 6767 14431 6792 14464
rect 6792 14431 6801 14464
rect 6839 14431 6860 14464
rect 6860 14431 6873 14464
rect 6911 14431 6928 14464
rect 6928 14431 6945 14464
rect 6983 14431 6996 14464
rect 6996 14431 7017 14464
rect 7055 14431 7064 14464
rect 7064 14431 7089 14464
rect 7127 14431 7132 14464
rect 7132 14431 7161 14464
rect 7199 14431 7200 14464
rect 7200 14431 7233 14464
rect 7271 14431 7302 14464
rect 7302 14431 7305 14464
rect 7343 14431 7370 14464
rect 7370 14431 7377 14464
rect 7415 14431 7438 14464
rect 7438 14431 7449 14464
rect 7487 14431 7506 14464
rect 7506 14431 7521 14464
rect 7559 14431 7574 14464
rect 7574 14431 7593 14464
rect 7631 14431 7642 14464
rect 7642 14431 7665 14464
rect 7703 14431 7710 14464
rect 7710 14431 7737 14464
rect 7775 14431 7778 14464
rect 7778 14431 7809 14464
rect 7847 14431 7880 14464
rect 7880 14431 7881 14464
rect 7919 14431 7948 14464
rect 7948 14431 7953 14464
rect 7991 14431 8016 14464
rect 8016 14431 8025 14464
rect 8063 14431 8084 14464
rect 8084 14431 8097 14464
rect 8135 14431 8152 14464
rect 8152 14431 8169 14464
rect 8207 14431 8220 14464
rect 8220 14431 8241 14464
rect 8279 14431 8288 14464
rect 8288 14431 8313 14464
rect 8351 14431 8356 14464
rect 8356 14431 8385 14464
rect 8423 14431 8424 14464
rect 8424 14431 8457 14464
rect 8495 14431 8526 14464
rect 8526 14431 8529 14464
rect 8567 14431 8594 14464
rect 8594 14431 8601 14464
rect 8639 14431 8662 14464
rect 8662 14431 8673 14464
rect 8711 14431 8730 14464
rect 8730 14431 8745 14464
rect 8783 14431 8798 14464
rect 8798 14431 8817 14464
rect 8855 14431 8866 14464
rect 8866 14431 8889 14464
rect 8927 14431 8934 14464
rect 8934 14431 8961 14464
rect 8999 14431 9002 14464
rect 9002 14431 9033 14464
rect 9071 14431 9104 14464
rect 9104 14431 9105 14464
rect 9143 14431 9172 14464
rect 9172 14431 9177 14464
rect 9215 14431 9240 14464
rect 9240 14431 9249 14464
rect 9287 14431 9308 14464
rect 9308 14431 9321 14464
rect 9359 14431 9376 14464
rect 9376 14431 9393 14464
rect 9431 14431 9444 14464
rect 9444 14431 9465 14464
rect 9503 14431 9512 14464
rect 9512 14431 9537 14464
rect 9575 14431 9580 14464
rect 9580 14431 9609 14464
rect 9647 14431 9648 14464
rect 9648 14431 9681 14464
rect 9719 14431 9750 14464
rect 9750 14431 9753 14464
rect 9791 14431 9818 14464
rect 9818 14431 9825 14464
rect 9863 14431 9886 14464
rect 9886 14431 9897 14464
rect 9935 14431 9954 14464
rect 9954 14431 9969 14464
rect 10007 14431 10022 14464
rect 10022 14431 10041 14464
rect 10079 14431 10090 14464
rect 10090 14431 10113 14464
rect 10151 14431 10158 14464
rect 10158 14431 10185 14464
rect 10223 14431 10226 14464
rect 10226 14431 10257 14464
rect 10295 14431 10328 14464
rect 10328 14431 10329 14464
rect 10367 14431 10396 14464
rect 10396 14431 10401 14464
rect 10439 14431 10464 14464
rect 10464 14431 10473 14464
rect 10511 14431 10532 14464
rect 10532 14431 10545 14464
rect 10583 14431 10600 14464
rect 10600 14431 10617 14464
rect 10655 14431 10668 14464
rect 10668 14431 10689 14464
rect 10727 14431 10736 14464
rect 10736 14431 10761 14464
rect 10799 14431 10804 14464
rect 10804 14431 10833 14464
rect 10871 14431 10872 14464
rect 10872 14431 10905 14464
rect 10943 14431 10974 14464
rect 10974 14431 10977 14464
rect 11015 14431 11042 14464
rect 11042 14431 11049 14464
rect 11087 14431 11110 14464
rect 11110 14431 11121 14464
rect 11159 14431 11178 14464
rect 11178 14431 11193 14464
rect 11231 14431 11246 14464
rect 11246 14431 11265 14464
rect 11303 14431 11314 14464
rect 11314 14431 11337 14464
rect 11375 14431 11382 14464
rect 11382 14431 11409 14464
rect 11447 14431 11450 14464
rect 11450 14431 11481 14464
rect 11519 14431 11552 14464
rect 11552 14431 11553 14464
rect 11591 14431 11620 14464
rect 11620 14431 11625 14464
rect 11663 14431 11688 14464
rect 11688 14431 11697 14464
rect 11735 14431 11756 14464
rect 11756 14431 11769 14464
rect 11807 14431 11824 14464
rect 11824 14431 11841 14464
rect 11879 14431 11892 14464
rect 11892 14431 11913 14464
rect 11951 14431 11960 14464
rect 11960 14431 11985 14464
rect 12023 14431 12028 14464
rect 12028 14431 12057 14464
rect 12095 14431 12096 14464
rect 12096 14431 12129 14464
rect 12167 14431 12198 14464
rect 12198 14431 12201 14464
rect 12239 14431 12266 14464
rect 12266 14431 12273 14464
rect 12311 14431 12334 14464
rect 12334 14431 12345 14464
rect 12383 14431 12402 14464
rect 12402 14431 12417 14464
rect 12455 14431 12470 14464
rect 12470 14431 12489 14464
rect 12527 14431 12538 14464
rect 12538 14431 12561 14464
rect 12599 14431 12606 14464
rect 12606 14431 12633 14464
rect 14306 14431 14340 14465
rect 14606 14431 14640 14465
<< metal1 >>
rect 877 37224 2226 37271
rect 877 36587 949 37224
rect 237 36547 949 36587
rect 237 36513 312 36547
rect 346 36513 949 36547
rect 237 36511 949 36513
rect 2153 36587 2226 37224
rect 12744 37221 14093 37275
rect 12744 36587 12813 37221
rect 2153 36511 12813 36587
rect 14017 36587 14093 37221
rect 14017 36546 14716 36587
rect 14017 36512 14606 36546
rect 14640 36512 14716 36546
rect 14017 36511 14716 36512
rect 237 36477 548 36511
rect 582 36477 620 36511
rect 654 36477 692 36511
rect 726 36477 764 36511
rect 798 36477 836 36511
rect 870 36477 908 36511
rect 942 36477 949 36511
rect 2166 36477 2204 36511
rect 2238 36477 2276 36511
rect 2310 36477 2348 36511
rect 2382 36477 2420 36511
rect 2454 36477 2492 36511
rect 2526 36477 2564 36511
rect 2598 36477 2636 36511
rect 2670 36477 2708 36511
rect 2742 36477 2780 36511
rect 2814 36477 2852 36511
rect 2886 36477 2924 36511
rect 2958 36477 2996 36511
rect 3030 36477 3068 36511
rect 3102 36477 3140 36511
rect 3174 36477 3212 36511
rect 3246 36477 3284 36511
rect 3318 36477 3356 36511
rect 3390 36477 3428 36511
rect 3462 36477 3500 36511
rect 3534 36477 3572 36511
rect 3606 36477 3644 36511
rect 3678 36477 3716 36511
rect 3750 36477 3788 36511
rect 3822 36477 3860 36511
rect 3894 36477 3932 36511
rect 3966 36477 4004 36511
rect 4038 36477 4076 36511
rect 4110 36477 4148 36511
rect 4182 36477 4220 36511
rect 4254 36477 4292 36511
rect 4326 36477 4364 36511
rect 4398 36477 4436 36511
rect 4470 36477 4508 36511
rect 4542 36477 4580 36511
rect 4614 36477 4652 36511
rect 4686 36477 4724 36511
rect 4758 36477 4796 36511
rect 4830 36477 4868 36511
rect 4902 36477 4940 36511
rect 4974 36477 5012 36511
rect 5046 36477 5084 36511
rect 5118 36477 5156 36511
rect 5190 36477 5228 36511
rect 5262 36477 5300 36511
rect 5334 36477 5372 36511
rect 5406 36477 5444 36511
rect 5478 36477 5516 36511
rect 5550 36477 5588 36511
rect 5622 36477 5660 36511
rect 5694 36477 5732 36511
rect 5766 36477 5804 36511
rect 5838 36477 5876 36511
rect 5910 36477 5948 36511
rect 5982 36477 6020 36511
rect 6054 36477 6092 36511
rect 6126 36477 6164 36511
rect 6198 36477 6236 36511
rect 6270 36477 6308 36511
rect 6342 36477 6380 36511
rect 6414 36477 6452 36511
rect 6486 36477 6524 36511
rect 6558 36477 6596 36511
rect 6630 36477 6668 36511
rect 6702 36477 6740 36511
rect 6774 36477 6812 36511
rect 6846 36477 6884 36511
rect 6918 36477 6956 36511
rect 6990 36477 7028 36511
rect 7062 36477 7100 36511
rect 7134 36477 7172 36511
rect 7206 36477 7244 36511
rect 7278 36477 7316 36511
rect 7350 36477 7388 36511
rect 7422 36477 7460 36511
rect 7494 36477 7532 36511
rect 7566 36477 7604 36511
rect 7638 36477 7676 36511
rect 7710 36477 7748 36511
rect 7782 36477 7820 36511
rect 7854 36477 7892 36511
rect 7926 36477 7964 36511
rect 7998 36477 8036 36511
rect 8070 36477 8108 36511
rect 8142 36477 8180 36511
rect 8214 36477 8252 36511
rect 8286 36477 8324 36511
rect 8358 36477 8396 36511
rect 8430 36477 8468 36511
rect 8502 36477 8540 36511
rect 8574 36477 8612 36511
rect 8646 36477 8684 36511
rect 8718 36477 8756 36511
rect 8790 36477 8828 36511
rect 8862 36477 8900 36511
rect 8934 36477 8972 36511
rect 9006 36477 9044 36511
rect 9078 36477 9116 36511
rect 9150 36477 9188 36511
rect 9222 36477 9260 36511
rect 9294 36477 9332 36511
rect 9366 36477 9404 36511
rect 9438 36477 9476 36511
rect 9510 36477 9548 36511
rect 9582 36477 9620 36511
rect 9654 36477 9692 36511
rect 9726 36477 9764 36511
rect 9798 36477 9836 36511
rect 9870 36477 9908 36511
rect 9942 36477 9980 36511
rect 10014 36477 10052 36511
rect 10086 36477 10124 36511
rect 10158 36477 10196 36511
rect 10230 36477 10268 36511
rect 10302 36477 10340 36511
rect 10374 36477 10412 36511
rect 10446 36477 10484 36511
rect 10518 36477 10556 36511
rect 10590 36477 10628 36511
rect 10662 36477 10700 36511
rect 10734 36477 10772 36511
rect 10806 36477 10844 36511
rect 10878 36477 10916 36511
rect 10950 36477 10988 36511
rect 11022 36477 11060 36511
rect 11094 36477 11132 36511
rect 11166 36477 11204 36511
rect 11238 36477 11276 36511
rect 11310 36477 11348 36511
rect 11382 36477 11420 36511
rect 11454 36477 11492 36511
rect 11526 36477 11564 36511
rect 11598 36477 11636 36511
rect 11670 36477 11708 36511
rect 11742 36477 11780 36511
rect 11814 36477 11852 36511
rect 11886 36477 11924 36511
rect 11958 36477 11996 36511
rect 12030 36477 12068 36511
rect 12102 36477 12140 36511
rect 12174 36477 12212 36511
rect 12246 36477 12284 36511
rect 12318 36477 12356 36511
rect 12390 36477 12428 36511
rect 12462 36477 12500 36511
rect 12534 36477 12572 36511
rect 12606 36477 12644 36511
rect 12678 36477 12716 36511
rect 12750 36477 12788 36511
rect 14046 36477 14084 36511
rect 14118 36477 14156 36511
rect 14190 36477 14228 36511
rect 14262 36477 14300 36511
rect 14334 36477 14372 36511
rect 14406 36477 14716 36511
rect 237 36475 949 36477
rect 237 36441 312 36475
rect 346 36468 949 36475
rect 2153 36468 12813 36477
rect 346 36465 12813 36468
rect 14017 36474 14716 36477
rect 14017 36465 14606 36474
rect 346 36441 14606 36465
rect 237 36440 14606 36441
rect 14640 36440 14716 36474
rect 237 36402 14716 36440
rect 237 36294 422 36402
rect 237 36260 312 36294
rect 346 36260 422 36294
rect 237 36222 422 36260
rect 237 36188 312 36222
rect 346 36188 422 36222
rect 237 36150 422 36188
rect 237 36116 312 36150
rect 346 36116 422 36150
rect 237 36078 422 36116
rect 237 36044 312 36078
rect 346 36044 422 36078
rect 14531 36291 14716 36402
rect 14531 36257 14606 36291
rect 14640 36257 14716 36291
rect 14531 36219 14716 36257
rect 14531 36185 14606 36219
rect 14640 36185 14716 36219
rect 14531 36147 14716 36185
rect 14531 36113 14606 36147
rect 14640 36113 14716 36147
rect 14531 36075 14716 36113
rect 237 36006 422 36044
rect 237 35972 312 36006
rect 346 35972 422 36006
rect 237 35934 422 35972
rect 237 35900 312 35934
rect 346 35900 422 35934
rect 237 35862 422 35900
rect 237 35828 312 35862
rect 346 35828 422 35862
rect 237 35790 422 35828
rect 237 35756 312 35790
rect 346 35756 422 35790
rect 237 35718 422 35756
rect 237 35684 312 35718
rect 346 35684 422 35718
rect 237 35646 422 35684
rect 237 35612 312 35646
rect 346 35612 422 35646
rect 237 35574 422 35612
rect 237 35540 312 35574
rect 346 35540 422 35574
rect 237 35502 422 35540
rect 237 35468 312 35502
rect 346 35468 422 35502
rect 237 35430 422 35468
rect 237 35396 312 35430
rect 346 35396 422 35430
rect 237 35358 422 35396
rect 237 35324 312 35358
rect 346 35324 422 35358
rect 237 35286 422 35324
rect 237 35252 312 35286
rect 346 35252 422 35286
rect 237 35214 422 35252
rect 237 35180 312 35214
rect 346 35180 422 35214
rect 237 35142 422 35180
rect 237 35108 312 35142
rect 346 35108 422 35142
rect 237 35070 422 35108
rect 237 35036 312 35070
rect 346 35036 422 35070
rect 237 34998 422 35036
rect 237 34964 312 34998
rect 346 34964 422 34998
rect 237 34926 422 34964
rect 237 34892 312 34926
rect 346 34892 422 34926
rect 237 34854 422 34892
rect 237 34820 312 34854
rect 346 34820 422 34854
rect 237 34782 422 34820
rect 237 34748 312 34782
rect 346 34748 422 34782
rect 237 34710 422 34748
rect 237 34676 312 34710
rect 346 34676 422 34710
rect 237 34638 422 34676
rect 237 34604 312 34638
rect 346 34604 422 34638
rect 237 34566 422 34604
rect 237 34532 312 34566
rect 346 34532 422 34566
rect 237 34494 422 34532
rect 237 34460 312 34494
rect 346 34460 422 34494
rect 237 34422 422 34460
rect 237 34388 312 34422
rect 346 34388 422 34422
rect 237 34350 422 34388
rect 237 34316 312 34350
rect 346 34316 422 34350
rect 237 34278 422 34316
rect 237 34244 312 34278
rect 346 34244 422 34278
rect 237 34206 422 34244
rect 237 34172 312 34206
rect 346 34172 422 34206
rect 237 34134 422 34172
rect 237 34100 312 34134
rect 346 34100 422 34134
rect 237 34062 422 34100
rect 237 34028 312 34062
rect 346 34028 422 34062
rect 237 33990 422 34028
rect 237 33956 312 33990
rect 346 33956 422 33990
rect 237 33918 422 33956
rect 237 33884 312 33918
rect 346 33884 422 33918
rect 237 33846 422 33884
rect 237 33812 312 33846
rect 346 33812 422 33846
rect 237 33774 422 33812
rect 237 33740 312 33774
rect 346 33740 422 33774
rect 237 33702 422 33740
rect 237 33668 312 33702
rect 346 33668 422 33702
rect 237 33630 422 33668
rect 237 33596 312 33630
rect 346 33596 422 33630
rect 237 33558 422 33596
rect 237 33524 312 33558
rect 346 33524 422 33558
rect 237 33486 422 33524
rect 237 33452 312 33486
rect 346 33452 422 33486
rect 237 33414 422 33452
rect 237 33380 312 33414
rect 346 33380 422 33414
rect 237 33342 422 33380
rect 237 33308 312 33342
rect 346 33308 422 33342
rect 237 33270 422 33308
rect 237 33236 312 33270
rect 346 33236 422 33270
rect 237 33198 422 33236
rect 237 33164 312 33198
rect 346 33164 422 33198
rect 237 33126 422 33164
rect 237 33092 312 33126
rect 346 33092 422 33126
rect 237 33054 422 33092
rect 237 33020 312 33054
rect 346 33020 422 33054
rect 237 32982 422 33020
rect 237 32948 312 32982
rect 346 32948 422 32982
rect 237 32910 422 32948
rect 237 32876 312 32910
rect 346 32876 422 32910
rect 237 32838 422 32876
rect 237 32804 312 32838
rect 346 32804 422 32838
rect 237 32766 422 32804
rect 237 32732 312 32766
rect 346 32732 422 32766
rect 237 32694 422 32732
rect 237 32660 312 32694
rect 346 32660 422 32694
rect 237 32622 422 32660
rect 237 32588 312 32622
rect 346 32588 422 32622
rect 237 32550 422 32588
rect 237 32516 312 32550
rect 346 32516 422 32550
rect 237 32478 422 32516
rect 237 32444 312 32478
rect 346 32444 422 32478
rect 237 32406 422 32444
rect 237 32372 312 32406
rect 346 32372 422 32406
rect 237 32334 422 32372
rect 237 32300 312 32334
rect 346 32300 422 32334
rect 237 32262 422 32300
rect 237 32228 312 32262
rect 346 32228 422 32262
rect 237 32190 422 32228
rect 237 32156 312 32190
rect 346 32156 422 32190
rect 237 32118 422 32156
rect 237 32084 312 32118
rect 346 32084 422 32118
rect 237 32046 422 32084
rect 237 32012 312 32046
rect 346 32012 422 32046
rect 237 31974 422 32012
rect 237 31940 312 31974
rect 346 31940 422 31974
rect 237 31902 422 31940
rect 237 31868 312 31902
rect 346 31868 422 31902
rect 237 31830 422 31868
rect 237 31796 312 31830
rect 346 31796 422 31830
rect 237 31758 422 31796
rect 237 31724 312 31758
rect 346 31724 422 31758
rect 237 31686 422 31724
rect 237 31652 312 31686
rect 346 31652 422 31686
rect 237 31614 422 31652
rect 237 31580 312 31614
rect 346 31580 422 31614
rect 237 31542 422 31580
rect 237 31508 312 31542
rect 346 31508 422 31542
rect 237 31470 422 31508
rect 237 31436 312 31470
rect 346 31436 422 31470
rect 237 31398 422 31436
rect 237 31364 312 31398
rect 346 31364 422 31398
rect 237 31326 422 31364
rect 237 31292 312 31326
rect 346 31292 422 31326
rect 237 31254 422 31292
rect 237 31220 312 31254
rect 346 31220 422 31254
rect 237 31182 422 31220
rect 237 31148 312 31182
rect 346 31148 422 31182
rect 237 31110 422 31148
rect 237 31076 312 31110
rect 346 31076 422 31110
rect 237 31038 422 31076
rect 237 31004 312 31038
rect 346 31004 422 31038
rect 237 30966 422 31004
rect 237 30932 312 30966
rect 346 30932 422 30966
rect 237 30894 422 30932
rect 237 30860 312 30894
rect 346 30860 422 30894
rect 237 30822 422 30860
rect 237 30788 312 30822
rect 346 30788 422 30822
rect 237 30750 422 30788
rect 237 30716 312 30750
rect 346 30716 422 30750
rect 237 30678 422 30716
rect 237 30644 312 30678
rect 346 30644 422 30678
rect 237 30606 422 30644
rect 237 30572 312 30606
rect 346 30572 422 30606
rect 237 30534 422 30572
rect 237 30500 312 30534
rect 346 30500 422 30534
rect 237 30462 422 30500
rect 237 30428 312 30462
rect 346 30428 422 30462
rect 237 30390 422 30428
rect 237 30356 312 30390
rect 346 30356 422 30390
rect 237 30318 422 30356
rect 237 30284 312 30318
rect 346 30284 422 30318
rect 237 30246 422 30284
rect 237 30212 312 30246
rect 346 30212 422 30246
rect 237 30174 422 30212
rect 237 30140 312 30174
rect 346 30140 422 30174
rect 237 30102 422 30140
rect 237 30068 312 30102
rect 346 30068 422 30102
rect 237 30030 422 30068
rect 237 29996 312 30030
rect 346 29996 422 30030
rect 237 29958 422 29996
rect 237 29924 312 29958
rect 346 29924 422 29958
rect 237 29886 422 29924
rect 237 29852 312 29886
rect 346 29852 422 29886
rect 237 29814 422 29852
rect 237 29780 312 29814
rect 346 29780 422 29814
rect 237 29742 422 29780
rect 237 29708 312 29742
rect 346 29708 422 29742
rect 237 29670 422 29708
rect 237 29636 312 29670
rect 346 29636 422 29670
rect 237 29598 422 29636
rect 237 29564 312 29598
rect 346 29564 422 29598
rect 237 29526 422 29564
rect 237 29492 312 29526
rect 346 29492 422 29526
rect 237 29454 422 29492
rect 237 29420 312 29454
rect 346 29420 422 29454
rect 237 29382 422 29420
rect 237 29348 312 29382
rect 346 29348 422 29382
rect 237 29310 422 29348
rect 237 29276 312 29310
rect 346 29276 422 29310
rect 237 29238 422 29276
rect 237 29204 312 29238
rect 346 29204 422 29238
rect 237 29166 422 29204
rect 237 29132 312 29166
rect 346 29132 422 29166
rect 237 29094 422 29132
rect 237 29060 312 29094
rect 346 29060 422 29094
rect 237 29022 422 29060
rect 237 28988 312 29022
rect 346 28988 422 29022
rect 237 28950 422 28988
rect 237 28916 312 28950
rect 346 28916 422 28950
rect 237 28878 422 28916
rect 237 28844 312 28878
rect 346 28844 422 28878
rect 237 28806 422 28844
rect 237 28772 312 28806
rect 346 28772 422 28806
rect 237 28734 422 28772
rect 237 28700 312 28734
rect 346 28700 422 28734
rect 237 28662 422 28700
rect 237 28628 312 28662
rect 346 28628 422 28662
rect 237 28590 422 28628
rect 237 28556 312 28590
rect 346 28556 422 28590
rect 237 28518 422 28556
rect 237 28484 312 28518
rect 346 28484 422 28518
rect 237 28446 422 28484
rect 237 28412 312 28446
rect 346 28412 422 28446
rect 237 28374 422 28412
rect 237 28340 312 28374
rect 346 28340 422 28374
rect 237 28302 422 28340
rect 237 28268 312 28302
rect 346 28268 422 28302
rect 237 28230 422 28268
rect 237 28196 312 28230
rect 346 28196 422 28230
rect 237 28158 422 28196
rect 237 28124 312 28158
rect 346 28124 422 28158
rect 237 28086 422 28124
rect 237 28052 312 28086
rect 346 28052 422 28086
rect 237 28014 422 28052
rect 237 27980 312 28014
rect 346 27980 422 28014
rect 237 27942 422 27980
rect 237 27908 312 27942
rect 346 27908 422 27942
rect 237 27870 422 27908
rect 237 27836 312 27870
rect 346 27836 422 27870
rect 237 27798 422 27836
rect 237 27764 312 27798
rect 346 27764 422 27798
rect 237 27726 422 27764
rect 237 27692 312 27726
rect 346 27692 422 27726
rect 237 27654 422 27692
rect 237 27620 312 27654
rect 346 27620 422 27654
rect 237 27582 422 27620
rect 237 27548 312 27582
rect 346 27548 422 27582
rect 237 27510 422 27548
rect 237 27476 312 27510
rect 346 27476 422 27510
rect 237 27438 422 27476
rect 237 27404 312 27438
rect 346 27404 422 27438
rect 237 27366 422 27404
rect 237 27332 312 27366
rect 346 27332 422 27366
rect 237 27294 422 27332
rect 237 27260 312 27294
rect 346 27260 422 27294
rect 237 27222 422 27260
rect 237 27188 312 27222
rect 346 27188 422 27222
rect 237 27150 422 27188
rect 237 27116 312 27150
rect 346 27116 422 27150
rect 237 27078 422 27116
rect 237 27044 312 27078
rect 346 27044 422 27078
rect 237 27006 422 27044
rect 237 26972 312 27006
rect 346 26972 422 27006
rect 237 26934 422 26972
rect 237 26900 312 26934
rect 346 26900 422 26934
rect 237 26862 422 26900
rect 237 26828 312 26862
rect 346 26828 422 26862
rect 237 26790 422 26828
rect 237 26756 312 26790
rect 346 26756 422 26790
rect 237 26718 422 26756
rect 237 26684 312 26718
rect 346 26684 422 26718
rect 237 26646 422 26684
rect 237 26612 312 26646
rect 346 26612 422 26646
rect 237 26574 422 26612
rect 237 26540 312 26574
rect 346 26540 422 26574
rect 237 26502 422 26540
rect 237 26468 312 26502
rect 346 26468 422 26502
rect 237 26430 422 26468
rect 237 26396 312 26430
rect 346 26396 422 26430
rect 237 26358 422 26396
rect 237 26324 312 26358
rect 346 26324 422 26358
rect 237 26286 422 26324
rect 237 26252 312 26286
rect 346 26252 422 26286
rect 237 26214 422 26252
rect 237 26180 312 26214
rect 346 26180 422 26214
rect 237 26142 422 26180
rect 237 26108 312 26142
rect 346 26108 422 26142
rect 237 26070 422 26108
rect 237 26036 312 26070
rect 346 26036 422 26070
rect 237 25998 422 26036
rect 237 25964 312 25998
rect 346 25964 422 25998
rect 237 25926 422 25964
rect 237 25892 312 25926
rect 346 25892 422 25926
rect 237 25854 422 25892
rect 237 25820 312 25854
rect 346 25820 422 25854
rect 237 25782 422 25820
rect 237 25748 312 25782
rect 346 25748 422 25782
rect 237 25710 422 25748
rect 237 25676 312 25710
rect 346 25676 422 25710
rect 237 25638 422 25676
rect 237 25604 312 25638
rect 346 25604 422 25638
rect 237 25566 422 25604
rect 237 25532 312 25566
rect 346 25532 422 25566
rect 237 25494 422 25532
rect 237 25460 312 25494
rect 346 25460 422 25494
rect 237 25422 422 25460
rect 237 25388 312 25422
rect 346 25388 422 25422
rect 237 25350 422 25388
rect 237 25316 312 25350
rect 346 25316 422 25350
rect 237 25278 422 25316
rect 237 25244 312 25278
rect 346 25244 422 25278
rect 237 25206 422 25244
rect 237 25172 312 25206
rect 346 25172 422 25206
rect 237 25134 422 25172
rect 237 25100 312 25134
rect 346 25100 422 25134
rect 237 25062 422 25100
rect 237 25028 312 25062
rect 346 25028 422 25062
rect 237 24990 422 25028
rect 237 24956 312 24990
rect 346 24956 422 24990
rect 237 24918 422 24956
rect 237 24884 312 24918
rect 346 24884 422 24918
rect 237 24846 422 24884
rect 237 24812 312 24846
rect 346 24812 422 24846
rect 237 24774 422 24812
rect 237 24740 312 24774
rect 346 24740 422 24774
rect 237 24702 422 24740
rect 237 24668 312 24702
rect 346 24668 422 24702
rect 237 24630 422 24668
rect 237 24596 312 24630
rect 346 24596 422 24630
rect 237 24558 422 24596
rect 237 24524 312 24558
rect 346 24524 422 24558
rect 237 24486 422 24524
rect 237 24452 312 24486
rect 346 24452 422 24486
rect 237 24414 422 24452
rect 237 24380 312 24414
rect 346 24380 422 24414
rect 237 24342 422 24380
rect 237 24308 312 24342
rect 346 24308 422 24342
rect 237 24270 422 24308
rect 237 24236 312 24270
rect 346 24236 422 24270
rect 237 24198 422 24236
rect 237 24164 312 24198
rect 346 24164 422 24198
rect 237 24126 422 24164
rect 237 24092 312 24126
rect 346 24092 422 24126
rect 237 24054 422 24092
rect 237 24020 312 24054
rect 346 24020 422 24054
rect 237 23982 422 24020
rect 237 23948 312 23982
rect 346 23948 422 23982
rect 237 23910 422 23948
rect 237 23876 312 23910
rect 346 23876 422 23910
rect 237 23838 422 23876
rect 237 23804 312 23838
rect 346 23804 422 23838
rect 237 23766 422 23804
rect 237 23732 312 23766
rect 346 23732 422 23766
rect 237 23694 422 23732
rect 237 23660 312 23694
rect 346 23660 422 23694
rect 237 23622 422 23660
rect 237 23588 312 23622
rect 346 23588 422 23622
rect 237 23550 422 23588
rect 237 23516 312 23550
rect 346 23516 422 23550
rect 237 23478 422 23516
rect 237 23444 312 23478
rect 346 23444 422 23478
rect 237 23406 422 23444
rect 237 23372 312 23406
rect 346 23372 422 23406
rect 237 23334 422 23372
rect 237 23300 312 23334
rect 346 23300 422 23334
rect 237 23262 422 23300
rect 237 23228 312 23262
rect 346 23228 422 23262
rect 237 23190 422 23228
rect 237 23156 312 23190
rect 346 23156 422 23190
rect 237 23118 422 23156
rect 237 23084 312 23118
rect 346 23084 422 23118
rect 237 23046 422 23084
rect 237 23012 312 23046
rect 346 23012 422 23046
rect 237 22974 422 23012
rect 237 22940 312 22974
rect 346 22940 422 22974
rect 237 22902 422 22940
rect 237 22868 312 22902
rect 346 22868 422 22902
rect 237 22830 422 22868
rect 237 22796 312 22830
rect 346 22796 422 22830
rect 237 22758 422 22796
rect 237 22724 312 22758
rect 346 22724 422 22758
rect 237 22686 422 22724
rect 237 22652 312 22686
rect 346 22652 422 22686
rect 237 22614 422 22652
rect 237 22580 312 22614
rect 346 22580 422 22614
rect 237 22542 422 22580
rect 237 22508 312 22542
rect 346 22508 422 22542
rect 237 22470 422 22508
rect 237 22436 312 22470
rect 346 22436 422 22470
rect 237 22398 422 22436
rect 237 22364 312 22398
rect 346 22364 422 22398
rect 237 22326 422 22364
rect 237 22292 312 22326
rect 346 22292 422 22326
rect 237 22254 422 22292
rect 237 22220 312 22254
rect 346 22220 422 22254
rect 237 22182 422 22220
rect 237 22148 312 22182
rect 346 22148 422 22182
rect 237 22110 422 22148
rect 237 22076 312 22110
rect 346 22076 422 22110
rect 237 22038 422 22076
rect 237 22004 312 22038
rect 346 22004 422 22038
rect 237 21966 422 22004
rect 237 21932 312 21966
rect 346 21932 422 21966
rect 237 21894 422 21932
rect 237 21860 312 21894
rect 346 21860 422 21894
rect 237 21822 422 21860
rect 237 21788 312 21822
rect 346 21788 422 21822
rect 237 21750 422 21788
rect 237 21716 312 21750
rect 346 21716 422 21750
rect 237 21678 422 21716
rect 237 21644 312 21678
rect 346 21644 422 21678
rect 237 21606 422 21644
rect 237 21572 312 21606
rect 346 21572 422 21606
rect 237 21534 422 21572
rect 237 21500 312 21534
rect 346 21500 422 21534
rect 237 21462 422 21500
rect 237 21428 312 21462
rect 346 21428 422 21462
rect 237 21390 422 21428
rect 237 21356 312 21390
rect 346 21356 422 21390
rect 237 21318 422 21356
rect 237 21284 312 21318
rect 346 21284 422 21318
rect 237 21246 422 21284
rect 237 21212 312 21246
rect 346 21212 422 21246
rect 237 21174 422 21212
rect 237 21140 312 21174
rect 346 21140 422 21174
rect 237 21102 422 21140
rect 237 21068 312 21102
rect 346 21068 422 21102
rect 237 21030 422 21068
rect 237 20996 312 21030
rect 346 20996 422 21030
rect 237 20958 422 20996
rect 237 20924 312 20958
rect 346 20924 422 20958
rect 237 20886 422 20924
rect 237 20852 312 20886
rect 346 20852 422 20886
rect 237 20814 422 20852
rect 237 20780 312 20814
rect 346 20780 422 20814
rect 237 20742 422 20780
rect 237 20708 312 20742
rect 346 20708 422 20742
rect 237 20670 422 20708
rect 237 20636 312 20670
rect 346 20636 422 20670
rect 237 20598 422 20636
rect 237 20564 312 20598
rect 346 20564 422 20598
rect 237 20526 422 20564
rect 237 20492 312 20526
rect 346 20492 422 20526
rect 237 20454 422 20492
rect 237 20420 312 20454
rect 346 20420 422 20454
rect 237 20382 422 20420
rect 237 20348 312 20382
rect 346 20348 422 20382
rect 237 20310 422 20348
rect 237 20276 312 20310
rect 346 20276 422 20310
rect 237 20238 422 20276
rect 237 20204 312 20238
rect 346 20204 422 20238
rect 237 20166 422 20204
rect 237 20132 312 20166
rect 346 20132 422 20166
rect 237 20094 422 20132
rect 237 20060 312 20094
rect 346 20060 422 20094
rect 237 20022 422 20060
rect 237 19988 312 20022
rect 346 19988 422 20022
rect 237 19950 422 19988
rect 237 19916 312 19950
rect 346 19916 422 19950
rect 237 19878 422 19916
rect 237 19844 312 19878
rect 346 19844 422 19878
rect 237 19806 422 19844
rect 237 19772 312 19806
rect 346 19772 422 19806
rect 237 19734 422 19772
rect 237 19700 312 19734
rect 346 19700 422 19734
rect 237 19662 422 19700
rect 237 19628 312 19662
rect 346 19628 422 19662
rect 237 19590 422 19628
rect 237 19556 312 19590
rect 346 19556 422 19590
rect 237 19518 422 19556
rect 237 19484 312 19518
rect 346 19484 422 19518
rect 237 19446 422 19484
rect 237 19412 312 19446
rect 346 19412 422 19446
rect 237 19374 422 19412
rect 237 19340 312 19374
rect 346 19340 422 19374
rect 237 19302 422 19340
rect 237 19268 312 19302
rect 346 19268 422 19302
rect 237 19230 422 19268
rect 237 19196 312 19230
rect 346 19196 422 19230
rect 237 19158 422 19196
rect 237 19124 312 19158
rect 346 19124 422 19158
rect 237 19086 422 19124
rect 237 19052 312 19086
rect 346 19052 422 19086
rect 237 19014 422 19052
rect 237 18980 312 19014
rect 346 18980 422 19014
rect 237 18942 422 18980
rect 237 18908 312 18942
rect 346 18908 422 18942
rect 237 18870 422 18908
rect 237 18836 312 18870
rect 346 18836 422 18870
rect 237 18798 422 18836
rect 237 18764 312 18798
rect 346 18764 422 18798
rect 237 18726 422 18764
rect 237 18692 312 18726
rect 346 18692 422 18726
rect 237 18654 422 18692
rect 237 18620 312 18654
rect 346 18620 422 18654
rect 237 18582 422 18620
rect 237 18548 312 18582
rect 346 18548 422 18582
rect 237 18510 422 18548
rect 237 18476 312 18510
rect 346 18476 422 18510
rect 237 18438 422 18476
rect 237 18404 312 18438
rect 346 18404 422 18438
rect 237 18366 422 18404
rect 237 18332 312 18366
rect 346 18332 422 18366
rect 237 18294 422 18332
rect 237 18260 312 18294
rect 346 18260 422 18294
rect 237 18222 422 18260
rect 237 18188 312 18222
rect 346 18188 422 18222
rect 237 18150 422 18188
rect 237 18116 312 18150
rect 346 18116 422 18150
rect 237 18078 422 18116
rect 237 18044 312 18078
rect 346 18044 422 18078
rect 237 18006 422 18044
rect 237 17972 312 18006
rect 346 17972 422 18006
rect 237 17934 422 17972
rect 237 17900 312 17934
rect 346 17900 422 17934
rect 237 17862 422 17900
rect 237 17828 312 17862
rect 346 17828 422 17862
rect 237 17790 422 17828
rect 237 17756 312 17790
rect 346 17756 422 17790
rect 237 17718 422 17756
rect 237 17684 312 17718
rect 346 17684 422 17718
rect 237 17646 422 17684
rect 237 17612 312 17646
rect 346 17612 422 17646
rect 237 17574 422 17612
rect 237 17540 312 17574
rect 346 17540 422 17574
rect 237 17502 422 17540
rect 237 17468 312 17502
rect 346 17468 422 17502
rect 237 17430 422 17468
rect 237 17396 312 17430
rect 346 17396 422 17430
rect 237 17358 422 17396
rect 237 17324 312 17358
rect 346 17324 422 17358
rect 237 17286 422 17324
rect 237 17252 312 17286
rect 346 17252 422 17286
rect 237 17214 422 17252
rect 237 17180 312 17214
rect 346 17180 422 17214
rect 237 17142 422 17180
rect 237 17108 312 17142
rect 346 17108 422 17142
rect 237 17070 422 17108
rect 237 17036 312 17070
rect 346 17036 422 17070
rect 237 16998 422 17036
rect 237 16964 312 16998
rect 346 16964 422 16998
rect 237 16926 422 16964
rect 237 16892 312 16926
rect 346 16892 422 16926
rect 237 16854 422 16892
rect 237 16820 312 16854
rect 346 16820 422 16854
rect 237 16782 422 16820
rect 237 16748 312 16782
rect 346 16748 422 16782
rect 237 16710 422 16748
rect 237 16676 312 16710
rect 346 16676 422 16710
rect 237 16638 422 16676
rect 237 16604 312 16638
rect 346 16604 422 16638
rect 237 16566 422 16604
rect 237 16532 312 16566
rect 346 16532 422 16566
rect 237 16494 422 16532
rect 237 16460 312 16494
rect 346 16460 422 16494
rect 237 16422 422 16460
rect 237 16388 312 16422
rect 346 16388 422 16422
rect 237 16350 422 16388
rect 237 16316 312 16350
rect 346 16316 422 16350
rect 237 16278 422 16316
rect 237 16244 312 16278
rect 346 16244 422 16278
rect 237 16206 422 16244
rect 237 16172 312 16206
rect 346 16172 422 16206
rect 237 16134 422 16172
rect 237 16100 312 16134
rect 346 16100 422 16134
rect 237 16062 422 16100
rect 237 16028 312 16062
rect 346 16028 422 16062
rect 237 15990 422 16028
rect 237 15956 312 15990
rect 346 15956 422 15990
rect 237 15918 422 15956
rect 237 15884 312 15918
rect 346 15884 422 15918
rect 237 15846 422 15884
rect 237 15812 312 15846
rect 346 15812 422 15846
rect 237 15774 422 15812
rect 237 15740 312 15774
rect 346 15740 422 15774
rect 237 15702 422 15740
rect 237 15668 312 15702
rect 346 15668 422 15702
rect 237 15630 422 15668
rect 237 15596 312 15630
rect 346 15596 422 15630
rect 237 15558 422 15596
rect 237 15524 312 15558
rect 346 15524 422 15558
rect 237 15486 422 15524
rect 237 15452 312 15486
rect 346 15452 422 15486
rect 237 15414 422 15452
rect 237 15380 312 15414
rect 346 15380 422 15414
rect 237 15342 422 15380
rect 237 15308 312 15342
rect 346 15308 422 15342
rect 237 15270 422 15308
rect 237 15236 312 15270
rect 346 15236 422 15270
rect 237 15198 422 15236
rect 237 15164 312 15198
rect 346 15164 422 15198
rect 237 15126 422 15164
rect 237 15092 312 15126
rect 346 15092 422 15126
rect 237 15054 422 15092
rect 237 15020 312 15054
rect 346 15020 422 15054
rect 237 14982 422 15020
rect 237 14948 312 14982
rect 346 14948 422 14982
rect 237 14910 422 14948
rect 237 14876 312 14910
rect 346 14876 422 14910
rect 237 14838 422 14876
tri 749 35966 849 36066 se
rect 849 36016 14111 36066
rect 849 35982 1001 36016
rect 1035 35982 1073 36016
rect 1107 35982 1145 36016
rect 1179 35982 1217 36016
rect 1251 35982 1289 36016
rect 1323 35982 1361 36016
rect 1395 35982 1433 36016
rect 1467 35982 1505 36016
rect 1539 35982 1577 36016
rect 1611 35982 1649 36016
rect 1683 35982 1721 36016
rect 1755 35982 1793 36016
rect 1827 35982 1865 36016
rect 1899 35982 1937 36016
rect 1971 35982 2009 36016
rect 2043 35982 2081 36016
rect 2115 35982 2153 36016
rect 2187 35982 2225 36016
rect 2259 35982 2297 36016
rect 2331 35982 2369 36016
rect 2403 35982 2441 36016
rect 2475 35982 2513 36016
rect 2547 35982 2585 36016
rect 2619 35982 2657 36016
rect 2691 35982 2729 36016
rect 2763 35982 2801 36016
rect 2835 35982 2873 36016
rect 2907 35982 2945 36016
rect 2979 35982 3017 36016
rect 3051 35982 3089 36016
rect 3123 35982 3161 36016
rect 3195 35982 3233 36016
rect 3267 35982 3305 36016
rect 3339 35982 3377 36016
rect 3411 35982 3449 36016
rect 3483 35982 3521 36016
rect 3555 35982 3593 36016
rect 3627 35982 3665 36016
rect 3699 35982 3737 36016
rect 3771 35982 3809 36016
rect 3843 35982 3881 36016
rect 3915 35982 3953 36016
rect 3987 35982 4025 36016
rect 4059 35982 4097 36016
rect 4131 35982 4169 36016
rect 4203 35982 4241 36016
rect 4275 35982 4313 36016
rect 4347 35982 4385 36016
rect 4419 35982 4457 36016
rect 4491 35982 4529 36016
rect 4563 35982 4601 36016
rect 4635 35982 4673 36016
rect 4707 35982 4745 36016
rect 4779 35982 4817 36016
rect 4851 35982 4889 36016
rect 4923 35982 4961 36016
rect 4995 35982 5033 36016
rect 5067 35982 5105 36016
rect 5139 35982 5177 36016
rect 5211 35982 5249 36016
rect 5283 35982 5321 36016
rect 5355 35982 5393 36016
rect 5427 35982 5465 36016
rect 5499 35982 5537 36016
rect 5571 35982 5609 36016
rect 5643 35982 5681 36016
rect 5715 35982 5753 36016
rect 5787 35982 5825 36016
rect 5859 35982 5897 36016
rect 5931 35982 5969 36016
rect 6003 35982 6041 36016
rect 6075 35982 6113 36016
rect 6147 35982 6185 36016
rect 6219 35982 6257 36016
rect 6291 35982 6329 36016
rect 6363 35982 6401 36016
rect 6435 35982 6473 36016
rect 6507 35982 6545 36016
rect 6579 35982 6617 36016
rect 6651 35982 6689 36016
rect 6723 35982 6761 36016
rect 6795 35982 6833 36016
rect 6867 35982 6905 36016
rect 6939 35982 6977 36016
rect 7011 35982 7049 36016
rect 7083 35982 7121 36016
rect 7155 35982 7193 36016
rect 7227 35982 7265 36016
rect 7299 35982 7337 36016
rect 7371 35982 7409 36016
rect 7443 35982 7481 36016
rect 7515 35982 7553 36016
rect 7587 35982 7625 36016
rect 7659 35982 7697 36016
rect 7731 35982 7769 36016
rect 7803 35982 7841 36016
rect 7875 35982 7913 36016
rect 7947 35982 7985 36016
rect 8019 35982 8057 36016
rect 8091 35982 8129 36016
rect 8163 35982 8201 36016
rect 8235 35982 8273 36016
rect 8307 35982 8345 36016
rect 8379 35982 8417 36016
rect 8451 35982 8489 36016
rect 8523 35982 8561 36016
rect 8595 35982 8633 36016
rect 8667 35982 8705 36016
rect 8739 35982 8777 36016
rect 8811 35982 8849 36016
rect 8883 35982 8921 36016
rect 8955 35982 8993 36016
rect 9027 35982 9065 36016
rect 9099 35982 9137 36016
rect 9171 35982 9209 36016
rect 9243 35982 9281 36016
rect 9315 35982 9353 36016
rect 9387 35982 9425 36016
rect 9459 35982 9497 36016
rect 9531 35982 9569 36016
rect 9603 35982 9641 36016
rect 9675 35982 9713 36016
rect 9747 35982 9785 36016
rect 9819 35982 9857 36016
rect 9891 35982 9929 36016
rect 9963 35982 10001 36016
rect 10035 35982 10073 36016
rect 10107 35982 10145 36016
rect 10179 35982 10217 36016
rect 10251 35982 10289 36016
rect 10323 35982 10361 36016
rect 10395 35982 10433 36016
rect 10467 35982 10505 36016
rect 10539 35982 10577 36016
rect 10611 35982 10649 36016
rect 10683 35982 10721 36016
rect 10755 35982 10793 36016
rect 10827 35982 10865 36016
rect 10899 35982 10937 36016
rect 10971 35982 11009 36016
rect 11043 35982 11081 36016
rect 11115 35982 11153 36016
rect 11187 35982 11225 36016
rect 11259 35982 11297 36016
rect 11331 35982 11369 36016
rect 11403 35982 11441 36016
rect 11475 35982 11513 36016
rect 11547 35982 11585 36016
rect 11619 35982 11657 36016
rect 11691 35982 11729 36016
rect 11763 35982 11801 36016
rect 11835 35982 11873 36016
rect 11907 35982 11945 36016
rect 11979 35982 12017 36016
rect 12051 35982 12089 36016
rect 12123 35982 12161 36016
rect 12195 35982 12233 36016
rect 12267 35982 12305 36016
rect 12339 35982 12377 36016
rect 12411 35982 12449 36016
rect 12483 35982 12521 36016
rect 12555 35982 12593 36016
rect 12627 35982 12665 36016
rect 12699 35982 12737 36016
rect 12771 35982 12809 36016
rect 12843 35982 12881 36016
rect 12915 35982 12953 36016
rect 12987 35982 13025 36016
rect 13059 35982 13097 36016
rect 13131 35982 13169 36016
rect 13203 35982 13241 36016
rect 13275 35982 13313 36016
rect 13347 35982 13385 36016
rect 13419 35982 13457 36016
rect 13491 35982 13529 36016
rect 13563 35982 13601 36016
rect 13635 35982 13673 36016
rect 13707 35982 13745 36016
rect 13779 35982 13817 36016
rect 13851 35982 13889 36016
rect 13923 35982 13961 36016
rect 13995 35982 14111 36016
rect 849 35966 14111 35982
tri 14111 35966 14211 36066 sw
rect 749 35946 14211 35966
rect 749 35913 869 35946
rect 749 35879 799 35913
rect 833 35879 869 35913
tri 869 35906 909 35946 nw
tri 14051 35906 14091 35946 ne
rect 749 35841 869 35879
rect 749 35807 799 35841
rect 833 35807 869 35841
rect 749 35769 869 35807
rect 749 35735 799 35769
rect 833 35735 869 35769
rect 749 35697 869 35735
rect 749 35663 799 35697
rect 833 35663 869 35697
rect 749 35625 869 35663
rect 749 35591 799 35625
rect 833 35591 869 35625
rect 749 35553 869 35591
rect 749 35519 799 35553
rect 833 35519 869 35553
rect 749 35481 869 35519
rect 749 35447 799 35481
rect 833 35447 869 35481
rect 749 35409 869 35447
rect 749 35375 799 35409
rect 833 35375 869 35409
rect 749 35337 869 35375
rect 749 35303 799 35337
rect 833 35303 869 35337
rect 749 35265 869 35303
rect 749 35231 799 35265
rect 833 35231 869 35265
rect 749 35193 869 35231
rect 749 35159 799 35193
rect 833 35159 869 35193
rect 749 35121 869 35159
rect 749 35087 799 35121
rect 833 35087 869 35121
rect 749 35049 869 35087
rect 749 35015 799 35049
rect 833 35015 869 35049
rect 749 34977 869 35015
rect 749 34943 799 34977
rect 833 34943 869 34977
rect 749 34905 869 34943
rect 749 34871 799 34905
rect 833 34871 869 34905
rect 749 34833 869 34871
rect 749 34799 799 34833
rect 833 34799 869 34833
rect 749 34761 869 34799
rect 749 34727 799 34761
rect 833 34727 869 34761
rect 14091 35834 14211 35946
rect 14091 35800 14114 35834
rect 14148 35800 14211 35834
rect 14091 35762 14211 35800
rect 14091 35728 14114 35762
rect 14148 35728 14211 35762
rect 14091 35690 14211 35728
rect 14091 35656 14114 35690
rect 14148 35656 14211 35690
rect 14091 35618 14211 35656
rect 14091 35584 14114 35618
rect 14148 35584 14211 35618
rect 14091 35546 14211 35584
rect 14091 35512 14114 35546
rect 14148 35512 14211 35546
rect 14091 35474 14211 35512
rect 14091 35440 14114 35474
rect 14148 35440 14211 35474
rect 14091 35402 14211 35440
rect 14091 35368 14114 35402
rect 14148 35368 14211 35402
rect 14091 35330 14211 35368
rect 14091 35296 14114 35330
rect 14148 35296 14211 35330
rect 14091 35258 14211 35296
rect 14091 35224 14114 35258
rect 14148 35224 14211 35258
rect 14091 35186 14211 35224
rect 14091 35152 14114 35186
rect 14148 35152 14211 35186
rect 14091 35114 14211 35152
rect 14091 35080 14114 35114
rect 14148 35080 14211 35114
rect 14091 35042 14211 35080
rect 14091 35008 14114 35042
rect 14148 35008 14211 35042
rect 14091 34970 14211 35008
rect 14091 34936 14114 34970
rect 14148 34936 14211 34970
rect 14091 34898 14211 34936
rect 14091 34864 14114 34898
rect 14148 34864 14211 34898
rect 14091 34826 14211 34864
rect 14091 34792 14114 34826
rect 14148 34792 14211 34826
rect 14091 34754 14211 34792
rect 749 34689 869 34727
rect 749 34655 799 34689
rect 833 34655 869 34689
rect 749 34617 869 34655
rect 749 34583 799 34617
rect 833 34583 869 34617
rect 749 34545 869 34583
rect 749 34511 799 34545
rect 833 34511 869 34545
rect 749 34473 869 34511
rect 749 34439 799 34473
rect 833 34439 869 34473
rect 749 34401 869 34439
rect 749 34367 799 34401
rect 833 34367 869 34401
rect 749 34329 869 34367
rect 749 34295 799 34329
rect 833 34295 869 34329
rect 749 34257 869 34295
rect 749 34223 799 34257
rect 833 34223 869 34257
rect 749 34185 869 34223
rect 749 34151 799 34185
rect 833 34151 869 34185
rect 749 34113 869 34151
rect 749 34079 799 34113
rect 833 34079 869 34113
rect 749 34041 869 34079
rect 749 34007 799 34041
rect 833 34007 869 34041
rect 749 33969 869 34007
rect 749 33935 799 33969
rect 833 33935 869 33969
rect 749 33897 869 33935
rect 749 33863 799 33897
rect 833 33863 869 33897
rect 749 33825 869 33863
rect 749 33791 799 33825
rect 833 33791 869 33825
rect 749 33753 869 33791
rect 749 33719 799 33753
rect 833 33719 869 33753
rect 749 33681 869 33719
rect 749 33647 799 33681
rect 833 33647 869 33681
rect 749 33609 869 33647
rect 749 33575 799 33609
rect 833 33575 869 33609
rect 749 33537 869 33575
rect 749 33503 799 33537
rect 833 33503 869 33537
rect 749 33465 869 33503
rect 749 33431 799 33465
rect 833 33431 869 33465
rect 749 33393 869 33431
rect 749 33359 799 33393
rect 833 33359 869 33393
rect 749 33321 869 33359
rect 749 33287 799 33321
rect 833 33287 869 33321
rect 749 33249 869 33287
rect 749 33215 799 33249
rect 833 33215 869 33249
rect 749 33177 869 33215
rect 749 33143 799 33177
rect 833 33143 869 33177
rect 749 33105 869 33143
rect 749 33071 799 33105
rect 833 33071 869 33105
rect 749 33033 869 33071
rect 749 32999 799 33033
rect 833 32999 869 33033
rect 749 32961 869 32999
rect 749 32927 799 32961
rect 833 32927 869 32961
rect 749 32889 869 32927
rect 749 32855 799 32889
rect 833 32855 869 32889
rect 749 32817 869 32855
rect 749 32783 799 32817
rect 833 32783 869 32817
rect 749 32745 869 32783
rect 749 32711 799 32745
rect 833 32711 869 32745
rect 749 32673 869 32711
rect 749 32639 799 32673
rect 833 32639 869 32673
rect 749 32601 869 32639
rect 749 32567 799 32601
rect 833 32567 869 32601
rect 749 32529 869 32567
rect 749 32495 799 32529
rect 833 32495 869 32529
rect 749 32457 869 32495
rect 749 32423 799 32457
rect 833 32423 869 32457
rect 749 32385 869 32423
rect 749 32351 799 32385
rect 833 32351 869 32385
rect 749 32313 869 32351
rect 749 32279 799 32313
rect 833 32279 869 32313
rect 749 32241 869 32279
rect 749 32207 799 32241
rect 833 32207 869 32241
rect 749 32169 869 32207
rect 749 32135 799 32169
rect 833 32135 869 32169
rect 749 32097 869 32135
rect 749 32063 799 32097
rect 833 32063 869 32097
rect 749 32025 869 32063
rect 749 31991 799 32025
rect 833 31991 869 32025
rect 749 31953 869 31991
rect 749 31919 799 31953
rect 833 31919 869 31953
rect 749 31881 869 31919
rect 749 31847 799 31881
rect 833 31847 869 31881
rect 749 31809 869 31847
rect 749 31775 799 31809
rect 833 31775 869 31809
rect 749 31737 869 31775
rect 749 31703 799 31737
rect 833 31703 869 31737
rect 749 31665 869 31703
rect 749 31631 799 31665
rect 833 31631 869 31665
rect 749 31593 869 31631
rect 749 31559 799 31593
rect 833 31559 869 31593
rect 749 31521 869 31559
rect 749 31487 799 31521
rect 833 31487 869 31521
rect 749 31449 869 31487
rect 749 31415 799 31449
rect 833 31415 869 31449
rect 749 31377 869 31415
rect 749 31343 799 31377
rect 833 31343 869 31377
rect 749 31305 869 31343
rect 749 31271 799 31305
rect 833 31271 869 31305
rect 749 31233 869 31271
rect 749 31199 799 31233
rect 833 31199 869 31233
rect 749 31161 869 31199
rect 749 31127 799 31161
rect 833 31127 869 31161
rect 749 31089 869 31127
rect 749 31055 799 31089
rect 833 31055 869 31089
rect 749 31017 869 31055
rect 749 30983 799 31017
rect 833 30983 869 31017
rect 749 30945 869 30983
rect 749 30911 799 30945
rect 833 30911 869 30945
rect 749 30873 869 30911
rect 749 30839 799 30873
rect 833 30839 869 30873
rect 749 30801 869 30839
rect 749 30767 799 30801
rect 833 30767 869 30801
rect 749 30729 869 30767
rect 749 30695 799 30729
rect 833 30695 869 30729
rect 749 30657 869 30695
rect 749 30623 799 30657
rect 833 30623 869 30657
rect 749 30585 869 30623
rect 749 30551 799 30585
rect 833 30551 869 30585
rect 749 30513 869 30551
rect 749 30479 799 30513
rect 833 30479 869 30513
rect 749 30441 869 30479
rect 749 30407 799 30441
rect 833 30407 869 30441
rect 749 30369 869 30407
rect 749 30335 799 30369
rect 833 30335 869 30369
rect 749 30297 869 30335
rect 749 30263 799 30297
rect 833 30263 869 30297
rect 749 30225 869 30263
rect 749 30191 799 30225
rect 833 30191 869 30225
rect 749 30153 869 30191
rect 749 30119 799 30153
rect 833 30119 869 30153
rect 749 30081 869 30119
rect 749 30047 799 30081
rect 833 30047 869 30081
rect 749 30009 869 30047
rect 749 29975 799 30009
rect 833 29975 869 30009
rect 749 29937 869 29975
rect 749 29903 799 29937
rect 833 29903 869 29937
rect 749 29865 869 29903
rect 749 29831 799 29865
rect 833 29831 869 29865
rect 749 29793 869 29831
rect 749 29759 799 29793
rect 833 29759 869 29793
rect 749 29721 869 29759
rect 749 29687 799 29721
rect 833 29687 869 29721
rect 749 29649 869 29687
rect 749 29615 799 29649
rect 833 29615 869 29649
rect 749 29577 869 29615
rect 749 29543 799 29577
rect 833 29543 869 29577
rect 749 29505 869 29543
rect 749 29471 799 29505
rect 833 29471 869 29505
rect 749 29433 869 29471
rect 749 29399 799 29433
rect 833 29399 869 29433
rect 749 29361 869 29399
rect 749 29327 799 29361
rect 833 29327 869 29361
rect 749 29289 869 29327
rect 749 29255 799 29289
rect 833 29255 869 29289
rect 749 29217 869 29255
rect 749 29183 799 29217
rect 833 29183 869 29217
rect 749 29145 869 29183
rect 749 29111 799 29145
rect 833 29111 869 29145
rect 749 29073 869 29111
rect 749 29039 799 29073
rect 833 29039 869 29073
rect 749 29001 869 29039
rect 749 28967 799 29001
rect 833 28967 869 29001
rect 749 28929 869 28967
rect 749 28895 799 28929
rect 833 28895 869 28929
rect 749 28857 869 28895
rect 749 28823 799 28857
rect 833 28823 869 28857
rect 749 28785 869 28823
rect 749 28751 799 28785
rect 833 28751 869 28785
rect 749 28713 869 28751
rect 749 28679 799 28713
rect 833 28679 869 28713
rect 749 28641 869 28679
rect 749 28607 799 28641
rect 833 28607 869 28641
rect 749 28569 869 28607
rect 749 28535 799 28569
rect 833 28535 869 28569
rect 749 28497 869 28535
rect 749 28463 799 28497
rect 833 28463 869 28497
rect 749 28425 869 28463
rect 749 28391 799 28425
rect 833 28391 869 28425
rect 749 28353 869 28391
rect 749 28319 799 28353
rect 833 28319 869 28353
rect 749 28281 869 28319
rect 749 28247 799 28281
rect 833 28247 869 28281
rect 749 28209 869 28247
rect 749 28175 799 28209
rect 833 28175 869 28209
rect 749 28137 869 28175
rect 749 28103 799 28137
rect 833 28103 869 28137
rect 749 28065 869 28103
rect 749 28031 799 28065
rect 833 28031 869 28065
rect 749 27993 869 28031
rect 749 27959 799 27993
rect 833 27959 869 27993
rect 749 27921 869 27959
rect 749 27887 799 27921
rect 833 27887 869 27921
rect 749 27849 869 27887
rect 749 27815 799 27849
rect 833 27815 869 27849
rect 749 27777 869 27815
rect 749 27743 799 27777
rect 833 27743 869 27777
rect 749 27705 869 27743
rect 749 27671 799 27705
rect 833 27671 869 27705
rect 749 27633 869 27671
rect 749 27599 799 27633
rect 833 27599 869 27633
rect 749 27561 869 27599
rect 749 27527 799 27561
rect 833 27527 869 27561
rect 749 27489 869 27527
rect 749 27455 799 27489
rect 833 27455 869 27489
rect 749 27417 869 27455
rect 749 27383 799 27417
rect 833 27383 869 27417
rect 749 27345 869 27383
rect 749 27311 799 27345
rect 833 27311 869 27345
rect 749 27273 869 27311
rect 749 27239 799 27273
rect 833 27239 869 27273
rect 749 27201 869 27239
rect 749 27167 799 27201
rect 833 27167 869 27201
rect 749 27129 869 27167
rect 749 27095 799 27129
rect 833 27095 869 27129
rect 749 27057 869 27095
rect 749 27023 799 27057
rect 833 27023 869 27057
rect 749 26985 869 27023
rect 749 26951 799 26985
rect 833 26951 869 26985
rect 749 26913 869 26951
rect 749 26879 799 26913
rect 833 26879 869 26913
rect 749 26841 869 26879
rect 749 26807 799 26841
rect 833 26807 869 26841
rect 749 26769 869 26807
rect 749 26735 799 26769
rect 833 26735 869 26769
rect 749 26697 869 26735
rect 749 26663 799 26697
rect 833 26663 869 26697
rect 749 26625 869 26663
rect 749 26591 799 26625
rect 833 26591 869 26625
rect 749 26553 869 26591
rect 749 26519 799 26553
rect 833 26519 869 26553
rect 749 26481 869 26519
rect 749 26447 799 26481
rect 833 26447 869 26481
rect 749 26409 869 26447
rect 749 26375 799 26409
rect 833 26375 869 26409
rect 749 26337 869 26375
rect 749 26303 799 26337
rect 833 26303 869 26337
rect 749 26265 869 26303
rect 749 26231 799 26265
rect 833 26231 869 26265
rect 749 26193 869 26231
rect 749 26159 799 26193
rect 833 26159 869 26193
rect 749 26121 869 26159
rect 749 26087 799 26121
rect 833 26087 869 26121
rect 749 26049 869 26087
rect 749 26015 799 26049
rect 833 26015 869 26049
rect 749 25977 869 26015
rect 749 25943 799 25977
rect 833 25943 869 25977
rect 749 25905 869 25943
rect 749 25871 799 25905
rect 833 25871 869 25905
rect 749 25833 869 25871
rect 749 25799 799 25833
rect 833 25799 869 25833
rect 749 25761 869 25799
rect 749 25727 799 25761
rect 833 25727 869 25761
rect 749 25689 869 25727
rect 749 25655 799 25689
rect 833 25655 869 25689
rect 749 25617 869 25655
rect 749 25583 799 25617
rect 833 25583 869 25617
rect 749 25545 869 25583
rect 749 25511 799 25545
rect 833 25511 869 25545
rect 749 25473 869 25511
rect 749 25439 799 25473
rect 833 25439 869 25473
rect 749 25401 869 25439
rect 749 25367 799 25401
rect 833 25367 869 25401
rect 749 25329 869 25367
rect 749 25295 799 25329
rect 833 25295 869 25329
rect 749 25257 869 25295
rect 749 25223 799 25257
rect 833 25223 869 25257
rect 749 25185 869 25223
rect 749 25151 799 25185
rect 833 25151 869 25185
rect 749 25113 869 25151
rect 749 25079 799 25113
rect 833 25079 869 25113
rect 749 25041 869 25079
rect 749 25007 799 25041
rect 833 25007 869 25041
rect 749 24969 869 25007
rect 749 24935 799 24969
rect 833 24935 869 24969
rect 749 24897 869 24935
rect 749 24863 799 24897
rect 833 24863 869 24897
rect 749 24825 869 24863
rect 749 24791 799 24825
rect 833 24791 869 24825
rect 749 24753 869 24791
rect 749 24719 799 24753
rect 833 24719 869 24753
rect 749 24681 869 24719
rect 749 24647 799 24681
rect 833 24647 869 24681
rect 749 24609 869 24647
rect 749 24575 799 24609
rect 833 24575 869 24609
rect 749 24537 869 24575
rect 749 24503 799 24537
rect 833 24503 869 24537
rect 749 24465 869 24503
rect 749 24431 799 24465
rect 833 24431 869 24465
rect 749 24393 869 24431
rect 749 24359 799 24393
rect 833 24359 869 24393
rect 749 24321 869 24359
rect 749 24287 799 24321
rect 833 24287 869 24321
rect 749 24249 869 24287
rect 749 24215 799 24249
rect 833 24215 869 24249
rect 749 24177 869 24215
rect 749 24143 799 24177
rect 833 24143 869 24177
rect 749 24105 869 24143
rect 749 24071 799 24105
rect 833 24071 869 24105
rect 749 24033 869 24071
rect 749 23999 799 24033
rect 833 23999 869 24033
rect 749 23961 869 23999
rect 749 23927 799 23961
rect 833 23927 869 23961
rect 749 23889 869 23927
rect 749 23855 799 23889
rect 833 23855 869 23889
rect 749 23817 869 23855
rect 749 23783 799 23817
rect 833 23783 869 23817
rect 749 23745 869 23783
rect 749 23711 799 23745
rect 833 23711 869 23745
rect 749 23673 869 23711
rect 749 23639 799 23673
rect 833 23639 869 23673
rect 749 23601 869 23639
rect 749 23567 799 23601
rect 833 23567 869 23601
rect 749 23529 869 23567
rect 749 23495 799 23529
rect 833 23495 869 23529
rect 749 23457 869 23495
rect 749 23423 799 23457
rect 833 23423 869 23457
rect 749 23385 869 23423
rect 749 23351 799 23385
rect 833 23351 869 23385
rect 749 23313 869 23351
rect 749 23279 799 23313
rect 833 23279 869 23313
rect 749 23241 869 23279
rect 749 23207 799 23241
rect 833 23207 869 23241
rect 749 23169 869 23207
rect 749 23135 799 23169
rect 833 23135 869 23169
rect 749 23097 869 23135
rect 749 23063 799 23097
rect 833 23063 869 23097
rect 749 23025 869 23063
rect 749 22991 799 23025
rect 833 22991 869 23025
rect 749 22953 869 22991
rect 749 22919 799 22953
rect 833 22919 869 22953
rect 749 22881 869 22919
rect 749 22847 799 22881
rect 833 22847 869 22881
rect 749 22809 869 22847
rect 749 22775 799 22809
rect 833 22775 869 22809
rect 749 22737 869 22775
rect 749 22703 799 22737
rect 833 22703 869 22737
rect 749 22665 869 22703
rect 749 22631 799 22665
rect 833 22631 869 22665
rect 749 22593 869 22631
rect 749 22559 799 22593
rect 833 22559 869 22593
rect 749 22521 869 22559
rect 749 22487 799 22521
rect 833 22487 869 22521
rect 749 22449 869 22487
rect 749 22415 799 22449
rect 833 22415 869 22449
rect 749 22377 869 22415
rect 749 22343 799 22377
rect 833 22343 869 22377
rect 749 22305 869 22343
rect 749 22271 799 22305
rect 833 22271 869 22305
rect 749 22233 869 22271
rect 749 22199 799 22233
rect 833 22199 869 22233
rect 749 22161 869 22199
rect 749 22127 799 22161
rect 833 22127 869 22161
rect 749 22089 869 22127
rect 749 22055 799 22089
rect 833 22055 869 22089
rect 749 22017 869 22055
rect 749 21983 799 22017
rect 833 21983 869 22017
rect 749 21945 869 21983
rect 749 21911 799 21945
rect 833 21911 869 21945
rect 749 21873 869 21911
rect 749 21839 799 21873
rect 833 21839 869 21873
rect 749 21801 869 21839
rect 749 21767 799 21801
rect 833 21767 869 21801
rect 749 21729 869 21767
rect 749 21695 799 21729
rect 833 21695 869 21729
rect 749 21657 869 21695
rect 749 21623 799 21657
rect 833 21623 869 21657
rect 749 21585 869 21623
rect 749 21551 799 21585
rect 833 21551 869 21585
rect 749 21513 869 21551
rect 749 21479 799 21513
rect 833 21479 869 21513
rect 749 21441 869 21479
rect 749 21407 799 21441
rect 833 21407 869 21441
rect 749 21369 869 21407
rect 749 21335 799 21369
rect 833 21335 869 21369
rect 749 21297 869 21335
rect 749 21263 799 21297
rect 833 21263 869 21297
rect 749 21225 869 21263
rect 749 21191 799 21225
rect 833 21191 869 21225
rect 749 21153 869 21191
rect 749 21119 799 21153
rect 833 21119 869 21153
rect 749 21081 869 21119
rect 749 21047 799 21081
rect 833 21047 869 21081
rect 749 21009 869 21047
rect 749 20975 799 21009
rect 833 20975 869 21009
rect 749 20937 869 20975
rect 749 20903 799 20937
rect 833 20903 869 20937
rect 749 20865 869 20903
rect 749 20831 799 20865
rect 833 20831 869 20865
rect 749 20793 869 20831
rect 749 20759 799 20793
rect 833 20759 869 20793
rect 749 20721 869 20759
rect 749 20687 799 20721
rect 833 20687 869 20721
rect 749 20649 869 20687
rect 749 20615 799 20649
rect 833 20615 869 20649
rect 749 20577 869 20615
rect 749 20543 799 20577
rect 833 20543 869 20577
rect 749 20505 869 20543
rect 749 20471 799 20505
rect 833 20471 869 20505
rect 749 20433 869 20471
rect 749 20399 799 20433
rect 833 20399 869 20433
rect 749 20361 869 20399
rect 749 20327 799 20361
rect 833 20327 869 20361
rect 749 20289 869 20327
rect 749 20255 799 20289
rect 833 20255 869 20289
rect 749 20217 869 20255
rect 749 20183 799 20217
rect 833 20183 869 20217
rect 749 20145 869 20183
rect 749 20111 799 20145
rect 833 20111 869 20145
rect 749 20073 869 20111
rect 749 20039 799 20073
rect 833 20039 869 20073
rect 749 20001 869 20039
rect 749 19967 799 20001
rect 833 19967 869 20001
rect 749 19929 869 19967
rect 749 19895 799 19929
rect 833 19895 869 19929
rect 749 19857 869 19895
rect 749 19823 799 19857
rect 833 19823 869 19857
rect 749 19785 869 19823
rect 749 19751 799 19785
rect 833 19751 869 19785
rect 749 19713 869 19751
rect 749 19679 799 19713
rect 833 19679 869 19713
rect 749 19641 869 19679
rect 749 19607 799 19641
rect 833 19607 869 19641
rect 749 19569 869 19607
rect 749 19535 799 19569
rect 833 19535 869 19569
rect 749 19497 869 19535
rect 749 19463 799 19497
rect 833 19463 869 19497
rect 749 19425 869 19463
rect 749 19391 799 19425
rect 833 19391 869 19425
rect 749 19353 869 19391
rect 749 19319 799 19353
rect 833 19319 869 19353
rect 749 19281 869 19319
rect 749 19247 799 19281
rect 833 19247 869 19281
rect 749 19209 869 19247
rect 749 19175 799 19209
rect 833 19175 869 19209
rect 749 19137 869 19175
rect 749 19103 799 19137
rect 833 19103 869 19137
rect 749 19065 869 19103
rect 749 19031 799 19065
rect 833 19031 869 19065
rect 749 18993 869 19031
rect 749 18959 799 18993
rect 833 18959 869 18993
rect 749 18921 869 18959
rect 749 18887 799 18921
rect 833 18887 869 18921
rect 749 18849 869 18887
rect 749 18815 799 18849
rect 833 18815 869 18849
rect 749 18777 869 18815
rect 749 18743 799 18777
rect 833 18743 869 18777
rect 749 18705 869 18743
rect 749 18671 799 18705
rect 833 18671 869 18705
rect 749 18633 869 18671
rect 749 18599 799 18633
rect 833 18599 869 18633
rect 749 18561 869 18599
rect 749 18527 799 18561
rect 833 18527 869 18561
rect 749 18489 869 18527
rect 749 18455 799 18489
rect 833 18455 869 18489
rect 749 18417 869 18455
rect 749 18383 799 18417
rect 833 18383 869 18417
rect 749 18345 869 18383
rect 749 18311 799 18345
rect 833 18311 869 18345
rect 749 18273 869 18311
rect 749 18239 799 18273
rect 833 18239 869 18273
rect 749 18201 869 18239
rect 749 18167 799 18201
rect 833 18167 869 18201
rect 749 18129 869 18167
rect 749 18095 799 18129
rect 833 18095 869 18129
rect 749 18057 869 18095
rect 749 18023 799 18057
rect 833 18023 869 18057
rect 749 17985 869 18023
rect 749 17951 799 17985
rect 833 17951 869 17985
rect 749 17913 869 17951
rect 749 17879 799 17913
rect 833 17879 869 17913
rect 749 17841 869 17879
rect 749 17807 799 17841
rect 833 17807 869 17841
rect 749 17769 869 17807
rect 749 17735 799 17769
rect 833 17735 869 17769
rect 749 17697 869 17735
rect 749 17663 799 17697
rect 833 17663 869 17697
rect 749 17625 869 17663
rect 749 17591 799 17625
rect 833 17591 869 17625
rect 749 17553 869 17591
rect 749 17519 799 17553
rect 833 17519 869 17553
rect 749 17481 869 17519
rect 749 17447 799 17481
rect 833 17447 869 17481
rect 749 17409 869 17447
rect 749 17375 799 17409
rect 833 17375 869 17409
rect 749 17337 869 17375
rect 749 17303 799 17337
rect 833 17303 869 17337
rect 749 17265 869 17303
rect 749 17231 799 17265
rect 833 17231 869 17265
rect 749 17193 869 17231
rect 749 17159 799 17193
rect 833 17159 869 17193
rect 749 17121 869 17159
rect 749 17087 799 17121
rect 833 17087 869 17121
rect 749 17049 869 17087
rect 749 17015 799 17049
rect 833 17015 869 17049
rect 749 16977 869 17015
rect 749 16943 799 16977
rect 833 16943 869 16977
rect 749 16905 869 16943
rect 749 16871 799 16905
rect 833 16871 869 16905
rect 749 16833 869 16871
rect 749 16799 799 16833
rect 833 16799 869 16833
rect 749 16761 869 16799
rect 749 16727 799 16761
rect 833 16727 869 16761
rect 749 16689 869 16727
rect 749 16655 799 16689
rect 833 16655 869 16689
rect 749 16617 869 16655
rect 749 16583 799 16617
rect 833 16583 869 16617
rect 749 16545 869 16583
rect 749 16511 799 16545
rect 833 16511 869 16545
rect 749 16473 869 16511
rect 749 16439 799 16473
rect 833 16439 869 16473
rect 749 16401 869 16439
rect 749 16367 799 16401
rect 833 16367 869 16401
rect 749 16329 869 16367
rect 749 16295 799 16329
rect 833 16295 869 16329
rect 749 16257 869 16295
rect 749 16223 799 16257
rect 833 16223 869 16257
rect 749 16185 869 16223
rect 749 16151 799 16185
rect 833 16151 869 16185
rect 749 16113 869 16151
rect 749 16079 799 16113
rect 833 16079 869 16113
rect 749 16041 869 16079
rect 749 16007 799 16041
rect 833 16007 869 16041
rect 749 15969 869 16007
rect 749 15935 799 15969
rect 833 15935 869 15969
rect 749 15897 869 15935
rect 749 15863 799 15897
rect 833 15863 869 15897
rect 749 15825 869 15863
rect 749 15791 799 15825
rect 833 15791 869 15825
rect 749 15753 869 15791
rect 749 15719 799 15753
rect 833 15719 869 15753
rect 749 15681 869 15719
rect 749 15647 799 15681
rect 833 15647 869 15681
rect 749 15609 869 15647
rect 749 15575 799 15609
rect 833 15575 869 15609
rect 749 15537 869 15575
rect 749 15503 799 15537
rect 833 15503 869 15537
rect 749 15465 869 15503
rect 749 15431 799 15465
rect 833 15431 869 15465
rect 749 15393 869 15431
rect 749 15359 799 15393
rect 833 15359 869 15393
rect 749 15321 869 15359
rect 749 15287 799 15321
rect 833 15287 869 15321
rect 749 15249 869 15287
rect 749 15215 799 15249
rect 833 15215 869 15249
rect 749 15177 869 15215
rect 1111 34692 13879 34734
rect 1111 34658 1293 34692
rect 1327 34658 1365 34692
rect 1399 34658 1437 34692
rect 1471 34658 1509 34692
rect 1543 34658 1581 34692
rect 1615 34658 1653 34692
rect 1687 34658 1725 34692
rect 1759 34658 1797 34692
rect 1831 34658 1869 34692
rect 1903 34658 1941 34692
rect 1975 34658 2013 34692
rect 2047 34658 2085 34692
rect 2119 34658 2157 34692
rect 2191 34658 2229 34692
rect 2263 34658 2301 34692
rect 2335 34658 2373 34692
rect 2407 34658 2445 34692
rect 2479 34658 2517 34692
rect 2551 34658 2589 34692
rect 2623 34658 2661 34692
rect 2695 34658 2733 34692
rect 2767 34658 2805 34692
rect 2839 34658 2877 34692
rect 2911 34658 2949 34692
rect 2983 34658 3021 34692
rect 3055 34658 3093 34692
rect 3127 34658 3165 34692
rect 3199 34658 3237 34692
rect 3271 34658 3309 34692
rect 3343 34658 3381 34692
rect 3415 34658 3453 34692
rect 3487 34658 3525 34692
rect 3559 34658 3597 34692
rect 3631 34658 3669 34692
rect 3703 34658 3741 34692
rect 3775 34658 3813 34692
rect 3847 34658 3885 34692
rect 3919 34658 3957 34692
rect 3991 34658 4029 34692
rect 4063 34658 4101 34692
rect 4135 34658 4173 34692
rect 4207 34658 4245 34692
rect 4279 34658 4317 34692
rect 4351 34658 4389 34692
rect 4423 34658 4461 34692
rect 4495 34658 4533 34692
rect 4567 34658 4605 34692
rect 4639 34658 4677 34692
rect 4711 34658 4749 34692
rect 4783 34658 4821 34692
rect 4855 34658 4893 34692
rect 4927 34658 4965 34692
rect 4999 34658 5037 34692
rect 5071 34658 5109 34692
rect 5143 34658 5181 34692
rect 5215 34658 5253 34692
rect 5287 34658 5325 34692
rect 5359 34658 5397 34692
rect 5431 34658 5469 34692
rect 5503 34658 5541 34692
rect 5575 34658 5613 34692
rect 5647 34658 5685 34692
rect 5719 34658 5757 34692
rect 5791 34658 5829 34692
rect 5863 34658 5901 34692
rect 5935 34658 5973 34692
rect 6007 34658 6045 34692
rect 6079 34658 6117 34692
rect 6151 34658 6189 34692
rect 6223 34658 6261 34692
rect 6295 34658 6333 34692
rect 6367 34658 6405 34692
rect 6439 34658 6477 34692
rect 6511 34658 6549 34692
rect 6583 34658 6621 34692
rect 6655 34658 6693 34692
rect 6727 34658 6765 34692
rect 6799 34658 6837 34692
rect 6871 34658 6909 34692
rect 6943 34658 6981 34692
rect 7015 34658 7053 34692
rect 7087 34658 7125 34692
rect 7159 34658 7197 34692
rect 7231 34658 7269 34692
rect 7303 34658 7341 34692
rect 7375 34658 7413 34692
rect 7447 34658 7485 34692
rect 7519 34658 7557 34692
rect 7591 34658 7629 34692
rect 7663 34658 7701 34692
rect 7735 34658 7773 34692
rect 7807 34658 7845 34692
rect 7879 34658 7917 34692
rect 7951 34658 7989 34692
rect 8023 34658 8061 34692
rect 8095 34658 8133 34692
rect 8167 34658 8205 34692
rect 8239 34658 8277 34692
rect 8311 34658 8349 34692
rect 8383 34658 8421 34692
rect 8455 34658 8493 34692
rect 8527 34658 8565 34692
rect 8599 34658 8637 34692
rect 8671 34658 8709 34692
rect 8743 34658 8781 34692
rect 8815 34658 8853 34692
rect 8887 34658 8925 34692
rect 8959 34658 8997 34692
rect 9031 34658 9069 34692
rect 9103 34658 9141 34692
rect 9175 34658 9213 34692
rect 9247 34658 9285 34692
rect 9319 34658 9357 34692
rect 9391 34658 9429 34692
rect 9463 34658 9501 34692
rect 9535 34658 9573 34692
rect 9607 34658 9645 34692
rect 9679 34658 9717 34692
rect 9751 34658 9789 34692
rect 9823 34658 9861 34692
rect 9895 34658 9933 34692
rect 9967 34658 10005 34692
rect 10039 34658 10077 34692
rect 10111 34658 10149 34692
rect 10183 34658 10221 34692
rect 10255 34658 10293 34692
rect 10327 34658 10365 34692
rect 10399 34658 10437 34692
rect 10471 34658 10509 34692
rect 10543 34658 10581 34692
rect 10615 34658 10653 34692
rect 10687 34658 10725 34692
rect 10759 34658 10797 34692
rect 10831 34658 10869 34692
rect 10903 34658 10941 34692
rect 10975 34658 11013 34692
rect 11047 34658 11085 34692
rect 11119 34658 11157 34692
rect 11191 34658 11229 34692
rect 11263 34658 11301 34692
rect 11335 34658 11373 34692
rect 11407 34658 11445 34692
rect 11479 34658 11517 34692
rect 11551 34658 11589 34692
rect 11623 34658 11661 34692
rect 11695 34658 11733 34692
rect 11767 34658 11805 34692
rect 11839 34658 11877 34692
rect 11911 34658 11949 34692
rect 11983 34658 12021 34692
rect 12055 34658 12093 34692
rect 12127 34658 12165 34692
rect 12199 34658 12237 34692
rect 12271 34658 12309 34692
rect 12343 34658 12381 34692
rect 12415 34658 12453 34692
rect 12487 34658 12525 34692
rect 12559 34658 12597 34692
rect 12631 34658 12669 34692
rect 12703 34658 12741 34692
rect 12775 34658 12813 34692
rect 12847 34658 12885 34692
rect 12919 34658 12957 34692
rect 12991 34658 13029 34692
rect 13063 34658 13101 34692
rect 13135 34658 13173 34692
rect 13207 34658 13245 34692
rect 13279 34658 13317 34692
rect 13351 34658 13389 34692
rect 13423 34658 13461 34692
rect 13495 34658 13533 34692
rect 13567 34658 13605 34692
rect 13639 34658 13677 34692
rect 13711 34658 13879 34692
rect 1111 34616 13879 34658
rect 1111 34495 1229 34616
rect 1111 34461 1153 34495
rect 1187 34461 1229 34495
rect 1111 34423 1229 34461
rect 1111 34389 1153 34423
rect 1187 34389 1229 34423
rect 1111 34351 1229 34389
rect 1111 34317 1153 34351
rect 1187 34317 1229 34351
rect 1111 34279 1229 34317
rect 1111 34245 1153 34279
rect 1187 34245 1229 34279
rect 1111 34207 1229 34245
rect 1111 34173 1153 34207
rect 1187 34173 1229 34207
rect 1111 34135 1229 34173
rect 1111 34101 1153 34135
rect 1187 34101 1229 34135
rect 1111 34063 1229 34101
rect 1111 34029 1153 34063
rect 1187 34029 1229 34063
rect 1111 33991 1229 34029
rect 1111 33957 1153 33991
rect 1187 33957 1229 33991
rect 1111 33919 1229 33957
rect 1111 33885 1153 33919
rect 1187 33885 1229 33919
rect 1111 33847 1229 33885
rect 1111 33813 1153 33847
rect 1187 33813 1229 33847
rect 1111 33775 1229 33813
rect 1111 33741 1153 33775
rect 1187 33741 1229 33775
rect 1111 33703 1229 33741
rect 1111 33669 1153 33703
rect 1187 33669 1229 33703
rect 1111 33631 1229 33669
rect 1111 33597 1153 33631
rect 1187 33597 1229 33631
rect 1111 33559 1229 33597
rect 1111 33525 1153 33559
rect 1187 33525 1229 33559
rect 1111 33487 1229 33525
rect 1111 33453 1153 33487
rect 1187 33453 1229 33487
rect 1111 33415 1229 33453
rect 1111 33381 1153 33415
rect 1187 33381 1229 33415
rect 1111 33343 1229 33381
rect 1111 33309 1153 33343
rect 1187 33309 1229 33343
rect 1111 33271 1229 33309
rect 1111 33237 1153 33271
rect 1187 33237 1229 33271
rect 1111 33199 1229 33237
rect 1111 33165 1153 33199
rect 1187 33165 1229 33199
rect 1111 33127 1229 33165
rect 1111 33093 1153 33127
rect 1187 33093 1229 33127
rect 1111 33055 1229 33093
rect 1111 33021 1153 33055
rect 1187 33021 1229 33055
rect 1111 32983 1229 33021
rect 1111 32949 1153 32983
rect 1187 32949 1229 32983
rect 1111 32911 1229 32949
rect 1111 32877 1153 32911
rect 1187 32877 1229 32911
rect 1111 32839 1229 32877
rect 1111 32805 1153 32839
rect 1187 32805 1229 32839
rect 1111 32767 1229 32805
rect 1111 32733 1153 32767
rect 1187 32733 1229 32767
rect 1111 32695 1229 32733
rect 1111 32661 1153 32695
rect 1187 32661 1229 32695
rect 1111 32623 1229 32661
rect 1111 32589 1153 32623
rect 1187 32589 1229 32623
rect 1111 32551 1229 32589
rect 1111 32517 1153 32551
rect 1187 32517 1229 32551
rect 1111 32479 1229 32517
rect 1111 32445 1153 32479
rect 1187 32445 1229 32479
rect 1111 32407 1229 32445
rect 1111 32373 1153 32407
rect 1187 32373 1229 32407
rect 1111 32335 1229 32373
rect 1111 32301 1153 32335
rect 1187 32301 1229 32335
rect 1111 32263 1229 32301
rect 1111 32229 1153 32263
rect 1187 32229 1229 32263
rect 1111 32191 1229 32229
rect 1111 32157 1153 32191
rect 1187 32157 1229 32191
rect 1111 32119 1229 32157
rect 1111 32085 1153 32119
rect 1187 32085 1229 32119
rect 1111 32047 1229 32085
rect 1111 32013 1153 32047
rect 1187 32013 1229 32047
rect 1111 31975 1229 32013
rect 1111 31941 1153 31975
rect 1187 31941 1229 31975
rect 1111 31903 1229 31941
rect 1111 31869 1153 31903
rect 1187 31869 1229 31903
rect 1111 31831 1229 31869
rect 1111 31797 1153 31831
rect 1187 31797 1229 31831
rect 1111 31759 1229 31797
rect 1111 31725 1153 31759
rect 1187 31725 1229 31759
rect 1111 31687 1229 31725
rect 1111 31653 1153 31687
rect 1187 31653 1229 31687
rect 1111 31615 1229 31653
rect 1111 31581 1153 31615
rect 1187 31581 1229 31615
rect 1111 31543 1229 31581
rect 1111 31509 1153 31543
rect 1187 31509 1229 31543
rect 1111 31471 1229 31509
rect 1111 31437 1153 31471
rect 1187 31437 1229 31471
rect 1111 31399 1229 31437
rect 1111 31365 1153 31399
rect 1187 31365 1229 31399
rect 1111 31327 1229 31365
rect 1111 31293 1153 31327
rect 1187 31293 1229 31327
rect 1111 31255 1229 31293
rect 1111 31221 1153 31255
rect 1187 31221 1229 31255
rect 1111 31183 1229 31221
rect 1111 31149 1153 31183
rect 1187 31149 1229 31183
rect 1111 31111 1229 31149
rect 1111 31077 1153 31111
rect 1187 31077 1229 31111
rect 1111 31039 1229 31077
rect 1111 31005 1153 31039
rect 1187 31005 1229 31039
rect 1111 30967 1229 31005
rect 1111 30933 1153 30967
rect 1187 30933 1229 30967
rect 1111 30895 1229 30933
rect 1111 30861 1153 30895
rect 1187 30861 1229 30895
rect 1111 30823 1229 30861
rect 1111 30789 1153 30823
rect 1187 30789 1229 30823
rect 1111 30751 1229 30789
rect 1111 30717 1153 30751
rect 1187 30717 1229 30751
rect 1111 30679 1229 30717
rect 1111 30645 1153 30679
rect 1187 30645 1229 30679
rect 1111 30607 1229 30645
rect 1111 30573 1153 30607
rect 1187 30573 1229 30607
rect 1111 30535 1229 30573
rect 1111 30501 1153 30535
rect 1187 30501 1229 30535
rect 1111 30463 1229 30501
rect 1111 30429 1153 30463
rect 1187 30429 1229 30463
rect 1111 30391 1229 30429
rect 1111 30357 1153 30391
rect 1187 30357 1229 30391
rect 1111 30319 1229 30357
rect 1111 30285 1153 30319
rect 1187 30294 1229 30319
rect 13761 34487 13879 34616
rect 13761 34453 13801 34487
rect 13835 34453 13879 34487
rect 13761 34415 13879 34453
rect 13761 34381 13801 34415
rect 13835 34381 13879 34415
rect 13761 34343 13879 34381
rect 13761 34309 13801 34343
rect 13835 34309 13879 34343
rect 13761 34271 13879 34309
rect 13761 34237 13801 34271
rect 13835 34237 13879 34271
rect 13761 34199 13879 34237
rect 13761 34165 13801 34199
rect 13835 34165 13879 34199
rect 13761 34127 13879 34165
rect 13761 34093 13801 34127
rect 13835 34093 13879 34127
rect 13761 34055 13879 34093
rect 13761 34021 13801 34055
rect 13835 34021 13879 34055
rect 13761 33983 13879 34021
rect 13761 33949 13801 33983
rect 13835 33949 13879 33983
rect 13761 33911 13879 33949
rect 13761 33877 13801 33911
rect 13835 33877 13879 33911
rect 13761 33839 13879 33877
rect 13761 33805 13801 33839
rect 13835 33805 13879 33839
rect 13761 33767 13879 33805
rect 13761 33733 13801 33767
rect 13835 33733 13879 33767
rect 13761 33695 13879 33733
rect 13761 33661 13801 33695
rect 13835 33661 13879 33695
rect 13761 33623 13879 33661
rect 13761 33589 13801 33623
rect 13835 33589 13879 33623
rect 13761 33551 13879 33589
rect 13761 33517 13801 33551
rect 13835 33517 13879 33551
rect 13761 33479 13879 33517
rect 13761 33445 13801 33479
rect 13835 33445 13879 33479
rect 13761 33407 13879 33445
rect 13761 33373 13801 33407
rect 13835 33373 13879 33407
rect 13761 33335 13879 33373
rect 13761 33301 13801 33335
rect 13835 33301 13879 33335
rect 13761 33263 13879 33301
rect 13761 33229 13801 33263
rect 13835 33229 13879 33263
rect 13761 33191 13879 33229
rect 13761 33157 13801 33191
rect 13835 33157 13879 33191
rect 13761 33119 13879 33157
rect 13761 33085 13801 33119
rect 13835 33085 13879 33119
rect 13761 33047 13879 33085
rect 13761 33013 13801 33047
rect 13835 33013 13879 33047
rect 13761 32975 13879 33013
rect 13761 32941 13801 32975
rect 13835 32941 13879 32975
rect 13761 32903 13879 32941
rect 13761 32869 13801 32903
rect 13835 32869 13879 32903
rect 13761 32831 13879 32869
rect 13761 32797 13801 32831
rect 13835 32797 13879 32831
rect 13761 32759 13879 32797
rect 13761 32725 13801 32759
rect 13835 32725 13879 32759
rect 13761 32687 13879 32725
rect 13761 32653 13801 32687
rect 13835 32653 13879 32687
rect 13761 32615 13879 32653
rect 13761 32581 13801 32615
rect 13835 32581 13879 32615
rect 13761 32543 13879 32581
rect 13761 32509 13801 32543
rect 13835 32509 13879 32543
rect 13761 32471 13879 32509
rect 13761 32437 13801 32471
rect 13835 32437 13879 32471
rect 13761 32399 13879 32437
rect 13761 32365 13801 32399
rect 13835 32365 13879 32399
rect 13761 32327 13879 32365
rect 13761 32293 13801 32327
rect 13835 32293 13879 32327
rect 13761 32255 13879 32293
rect 13761 32221 13801 32255
rect 13835 32221 13879 32255
rect 13761 32183 13879 32221
rect 13761 32149 13801 32183
rect 13835 32149 13879 32183
rect 13761 32111 13879 32149
rect 13761 32077 13801 32111
rect 13835 32077 13879 32111
rect 13761 32039 13879 32077
rect 13761 32005 13801 32039
rect 13835 32005 13879 32039
rect 13761 31967 13879 32005
rect 13761 31933 13801 31967
rect 13835 31933 13879 31967
rect 13761 31895 13879 31933
rect 13761 31861 13801 31895
rect 13835 31861 13879 31895
rect 13761 31823 13879 31861
rect 13761 31789 13801 31823
rect 13835 31789 13879 31823
rect 13761 31751 13879 31789
rect 13761 31717 13801 31751
rect 13835 31717 13879 31751
rect 13761 31679 13879 31717
rect 13761 31645 13801 31679
rect 13835 31645 13879 31679
rect 13761 31607 13879 31645
rect 13761 31573 13801 31607
rect 13835 31573 13879 31607
rect 13761 31535 13879 31573
rect 13761 31501 13801 31535
rect 13835 31501 13879 31535
rect 13761 31463 13879 31501
rect 13761 31429 13801 31463
rect 13835 31429 13879 31463
rect 13761 31391 13879 31429
rect 13761 31357 13801 31391
rect 13835 31357 13879 31391
rect 13761 31319 13879 31357
rect 13761 31285 13801 31319
rect 13835 31285 13879 31319
rect 13761 31247 13879 31285
rect 13761 31213 13801 31247
rect 13835 31213 13879 31247
rect 13761 31175 13879 31213
rect 13761 31141 13801 31175
rect 13835 31141 13879 31175
rect 13761 31103 13879 31141
rect 13761 31069 13801 31103
rect 13835 31069 13879 31103
rect 13761 31031 13879 31069
rect 13761 30997 13801 31031
rect 13835 30997 13879 31031
rect 13761 30959 13879 30997
rect 13761 30925 13801 30959
rect 13835 30925 13879 30959
rect 13761 30887 13879 30925
rect 13761 30853 13801 30887
rect 13835 30853 13879 30887
rect 13761 30815 13879 30853
rect 13761 30781 13801 30815
rect 13835 30781 13879 30815
rect 13761 30743 13879 30781
rect 13761 30709 13801 30743
rect 13835 30709 13879 30743
rect 13761 30671 13879 30709
rect 13761 30637 13801 30671
rect 13835 30637 13879 30671
rect 13761 30599 13879 30637
rect 13761 30565 13801 30599
rect 13835 30565 13879 30599
rect 13761 30527 13879 30565
rect 13761 30493 13801 30527
rect 13835 30493 13879 30527
rect 13761 30455 13879 30493
rect 13761 30421 13801 30455
rect 13835 30421 13879 30455
rect 13761 30383 13879 30421
rect 13761 30349 13801 30383
rect 13835 30349 13879 30383
rect 13761 30311 13879 30349
rect 1187 30285 10083 30294
rect 1111 30247 10083 30285
rect 1111 30213 1153 30247
rect 1187 30240 10083 30247
rect 1187 30213 4936 30240
rect 1111 30175 4936 30213
rect 1111 30141 1153 30175
rect 1187 30141 4936 30175
rect 1111 30103 4936 30141
rect 1111 30069 1153 30103
rect 1187 30069 4936 30103
rect 1111 30031 4936 30069
rect 1111 29997 1153 30031
rect 1187 29997 4936 30031
rect 1111 29959 4936 29997
rect 1111 29925 1153 29959
rect 1187 29925 4936 29959
rect 1111 29887 4936 29925
rect 1111 29853 1153 29887
rect 1187 29853 4936 29887
rect 1111 29815 4936 29853
rect 1111 29781 1153 29815
rect 1187 29781 4936 29815
rect 1111 29743 4936 29781
rect 1111 29709 1153 29743
rect 1187 29709 4936 29743
rect 1111 29671 4936 29709
rect 1111 29637 1153 29671
rect 1187 29637 4936 29671
rect 1111 29599 4936 29637
rect 1111 29565 1153 29599
rect 1187 29565 4936 29599
rect 1111 29527 4936 29565
rect 1111 29493 1153 29527
rect 1187 29493 4936 29527
rect 1111 29455 4936 29493
rect 1111 29421 1153 29455
rect 1187 29421 4936 29455
rect 1111 29420 4936 29421
rect 7228 29420 7737 30240
rect 10029 30094 10083 30240
tri 10083 30094 10283 30294 sw
rect 10029 29566 10283 30094
rect 10029 29420 10083 29566
rect 1111 29383 10083 29420
rect 1111 29349 1153 29383
rect 1187 29366 10083 29383
tri 10083 29366 10283 29566 nw
rect 13761 30277 13801 30311
rect 13835 30277 13879 30311
rect 13761 30239 13879 30277
rect 13761 30205 13801 30239
rect 13835 30205 13879 30239
rect 13761 30167 13879 30205
rect 13761 30133 13801 30167
rect 13835 30133 13879 30167
rect 13761 30095 13879 30133
rect 13761 30061 13801 30095
rect 13835 30061 13879 30095
rect 13761 30023 13879 30061
rect 13761 29989 13801 30023
rect 13835 29989 13879 30023
rect 13761 29951 13879 29989
rect 13761 29917 13801 29951
rect 13835 29917 13879 29951
rect 13761 29879 13879 29917
rect 13761 29845 13801 29879
rect 13835 29845 13879 29879
rect 13761 29807 13879 29845
rect 13761 29773 13801 29807
rect 13835 29773 13879 29807
rect 13761 29735 13879 29773
rect 13761 29701 13801 29735
rect 13835 29701 13879 29735
rect 13761 29663 13879 29701
rect 13761 29629 13801 29663
rect 13835 29629 13879 29663
rect 13761 29591 13879 29629
rect 13761 29557 13801 29591
rect 13835 29557 13879 29591
rect 13761 29519 13879 29557
rect 13761 29485 13801 29519
rect 13835 29485 13879 29519
rect 13761 29447 13879 29485
rect 13761 29413 13801 29447
rect 13835 29413 13879 29447
rect 13761 29375 13879 29413
rect 1187 29349 1434 29366
rect 1111 29311 1434 29349
rect 1111 29277 1153 29311
rect 1187 29277 1434 29311
rect 1111 29239 1434 29277
rect 1111 29205 1153 29239
rect 1187 29205 1434 29239
rect 1111 29167 1434 29205
rect 1111 29133 1153 29167
rect 1187 29133 1434 29167
rect 1111 29095 1434 29133
rect 1111 29061 1153 29095
rect 1187 29061 1434 29095
rect 1111 29023 1434 29061
rect 1111 28989 1153 29023
rect 1187 28989 1434 29023
rect 1111 28951 1434 28989
rect 1111 28917 1153 28951
rect 1187 28917 1434 28951
rect 13761 29341 13801 29375
rect 13835 29341 13879 29375
rect 13761 29303 13879 29341
rect 13761 29269 13801 29303
rect 13835 29269 13879 29303
rect 13761 29231 13879 29269
rect 13761 29197 13801 29231
rect 13835 29197 13879 29231
rect 13761 29159 13879 29197
rect 13761 29125 13801 29159
rect 13835 29125 13879 29159
rect 13761 29087 13879 29125
rect 13761 29053 13801 29087
rect 13835 29053 13879 29087
rect 13761 29015 13879 29053
rect 13761 28981 13801 29015
rect 13835 28981 13879 29015
rect 13761 28943 13879 28981
rect 1111 28879 1434 28917
rect 1111 28845 1153 28879
rect 1187 28845 1434 28879
rect 1111 28807 1434 28845
rect 1111 28773 1153 28807
rect 1187 28773 1434 28807
rect 1111 28735 1434 28773
rect 1111 28701 1153 28735
rect 1187 28701 1434 28735
rect 1111 28663 1434 28701
rect 1111 28629 1153 28663
rect 1187 28629 1434 28663
rect 1111 28591 1434 28629
rect 1111 28557 1153 28591
rect 1187 28557 1434 28591
rect 1111 28519 1434 28557
rect 1111 28485 1153 28519
rect 1187 28485 1434 28519
rect 1111 28447 1434 28485
rect 1111 28413 1153 28447
rect 1187 28413 1434 28447
rect 1111 28375 1434 28413
rect 1111 28341 1153 28375
rect 1187 28341 1434 28375
rect 1111 28303 1434 28341
rect 1111 28269 1153 28303
rect 1187 28269 1434 28303
rect 1111 28231 1434 28269
rect 1111 28197 1153 28231
rect 1187 28197 1434 28231
rect 1111 28159 1434 28197
rect 1111 28125 1153 28159
rect 1187 28125 1434 28159
rect 1111 28087 1434 28125
rect 1111 28053 1153 28087
rect 1187 28053 1434 28087
rect 1111 28015 1434 28053
rect 1111 27981 1153 28015
rect 1187 27981 1434 28015
rect 1111 27943 1434 27981
rect 1111 27909 1153 27943
rect 1187 27909 1434 27943
rect 1111 27871 1434 27909
rect 1111 27837 1153 27871
rect 1187 27837 1434 27871
rect 1111 27799 1434 27837
rect 1111 27765 1153 27799
rect 1187 27765 1434 27799
rect 1111 27727 1434 27765
rect 1111 27693 1153 27727
rect 1187 27693 1434 27727
rect 1111 27655 1434 27693
rect 1111 27621 1153 27655
rect 1187 27621 1434 27655
rect 1111 27583 1434 27621
rect 1111 27549 1153 27583
rect 1187 27549 1434 27583
rect 1111 27511 1434 27549
rect 1111 27477 1153 27511
rect 1187 27477 1434 27511
rect 1111 27439 1434 27477
rect 1111 27405 1153 27439
rect 1187 27405 1434 27439
rect 1111 27367 1434 27405
rect 1111 27333 1153 27367
rect 1187 27333 1434 27367
rect 1111 27295 1434 27333
rect 1111 27261 1153 27295
rect 1187 27261 1434 27295
rect 1111 27223 1434 27261
rect 1111 27189 1153 27223
rect 1187 27189 1434 27223
rect 1111 27151 1434 27189
rect 1111 27117 1153 27151
rect 1187 27117 1434 27151
rect 1111 27079 1434 27117
rect 1111 27045 1153 27079
rect 1187 27045 1434 27079
rect 1111 27007 1434 27045
tri 1651 28722 1851 28922 se
rect 1851 28888 13149 28922
rect 1851 28722 1974 28888
rect 1651 28566 1974 28722
rect 13024 28566 13149 28888
rect 1651 28528 13149 28566
rect 1651 28502 2085 28528
rect 1651 27460 1718 28502
rect 1968 27460 2085 28502
tri 2085 28488 2125 28528 nw
tri 12875 28488 12915 28528 ne
rect 12915 28515 13149 28528
tri 13149 28515 13556 28922 sw
rect 13761 28909 13801 28943
rect 13835 28909 13879 28943
rect 13761 28871 13879 28909
rect 13761 28837 13801 28871
rect 13835 28837 13879 28871
rect 13761 28799 13879 28837
rect 13761 28765 13801 28799
rect 13835 28765 13879 28799
rect 13761 28740 13879 28765
rect 14091 34720 14114 34754
rect 14148 34720 14211 34754
rect 14091 34682 14211 34720
rect 14091 34648 14114 34682
rect 14148 34648 14211 34682
rect 14091 34610 14211 34648
rect 14091 34576 14114 34610
rect 14148 34576 14211 34610
rect 14091 34538 14211 34576
rect 14091 34504 14114 34538
rect 14148 34504 14211 34538
rect 14091 34466 14211 34504
rect 14091 34432 14114 34466
rect 14148 34432 14211 34466
rect 14091 34394 14211 34432
rect 14091 34360 14114 34394
rect 14148 34360 14211 34394
rect 14091 34322 14211 34360
rect 14091 34288 14114 34322
rect 14148 34288 14211 34322
rect 14091 34250 14211 34288
rect 14091 34216 14114 34250
rect 14148 34216 14211 34250
rect 14091 34178 14211 34216
rect 14091 34144 14114 34178
rect 14148 34144 14211 34178
rect 14091 34106 14211 34144
rect 14091 34072 14114 34106
rect 14148 34072 14211 34106
rect 14091 34034 14211 34072
rect 14091 34000 14114 34034
rect 14148 34000 14211 34034
rect 14091 33962 14211 34000
rect 14091 33928 14114 33962
rect 14148 33928 14211 33962
rect 14091 33890 14211 33928
rect 14091 33856 14114 33890
rect 14148 33856 14211 33890
rect 14091 33818 14211 33856
rect 14091 33784 14114 33818
rect 14148 33784 14211 33818
rect 14091 33746 14211 33784
rect 14091 33712 14114 33746
rect 14148 33712 14211 33746
rect 14091 33674 14211 33712
rect 14091 33640 14114 33674
rect 14148 33640 14211 33674
rect 14091 33602 14211 33640
rect 14091 33568 14114 33602
rect 14148 33568 14211 33602
rect 14091 33530 14211 33568
rect 14091 33496 14114 33530
rect 14148 33496 14211 33530
rect 14091 33458 14211 33496
rect 14091 33424 14114 33458
rect 14148 33424 14211 33458
rect 14091 33386 14211 33424
rect 14091 33352 14114 33386
rect 14148 33352 14211 33386
rect 14091 33314 14211 33352
rect 14091 33280 14114 33314
rect 14148 33280 14211 33314
rect 14091 33242 14211 33280
rect 14091 33208 14114 33242
rect 14148 33208 14211 33242
rect 14091 33170 14211 33208
rect 14091 33136 14114 33170
rect 14148 33136 14211 33170
rect 14091 33098 14211 33136
rect 14091 33064 14114 33098
rect 14148 33064 14211 33098
rect 14091 33026 14211 33064
rect 14091 32992 14114 33026
rect 14148 32992 14211 33026
rect 14091 32954 14211 32992
rect 14091 32920 14114 32954
rect 14148 32920 14211 32954
rect 14091 32882 14211 32920
rect 14091 32848 14114 32882
rect 14148 32848 14211 32882
rect 14091 32810 14211 32848
rect 14091 32776 14114 32810
rect 14148 32776 14211 32810
rect 14091 32738 14211 32776
rect 14091 32704 14114 32738
rect 14148 32704 14211 32738
rect 14091 32666 14211 32704
rect 14091 32632 14114 32666
rect 14148 32632 14211 32666
rect 14091 32594 14211 32632
rect 14091 32560 14114 32594
rect 14148 32560 14211 32594
rect 14091 32522 14211 32560
rect 14091 32488 14114 32522
rect 14148 32488 14211 32522
rect 14091 32450 14211 32488
rect 14091 32416 14114 32450
rect 14148 32416 14211 32450
rect 14091 32378 14211 32416
rect 14091 32344 14114 32378
rect 14148 32344 14211 32378
rect 14091 32306 14211 32344
rect 14091 32272 14114 32306
rect 14148 32272 14211 32306
rect 14091 32234 14211 32272
rect 14091 32200 14114 32234
rect 14148 32200 14211 32234
rect 14091 32162 14211 32200
rect 14091 32128 14114 32162
rect 14148 32128 14211 32162
rect 14091 32090 14211 32128
rect 14091 32056 14114 32090
rect 14148 32056 14211 32090
rect 14091 32018 14211 32056
rect 14091 31984 14114 32018
rect 14148 31984 14211 32018
rect 14091 31946 14211 31984
rect 14091 31912 14114 31946
rect 14148 31912 14211 31946
rect 14091 31874 14211 31912
rect 14091 31840 14114 31874
rect 14148 31840 14211 31874
rect 14091 31802 14211 31840
rect 14091 31768 14114 31802
rect 14148 31768 14211 31802
rect 14091 31730 14211 31768
rect 14091 31696 14114 31730
rect 14148 31696 14211 31730
rect 14091 31658 14211 31696
rect 14091 31624 14114 31658
rect 14148 31624 14211 31658
rect 14091 31586 14211 31624
rect 14091 31552 14114 31586
rect 14148 31552 14211 31586
rect 14091 31514 14211 31552
rect 14091 31480 14114 31514
rect 14148 31480 14211 31514
rect 14091 31442 14211 31480
rect 14091 31408 14114 31442
rect 14148 31408 14211 31442
rect 14091 31370 14211 31408
rect 14091 31336 14114 31370
rect 14148 31336 14211 31370
rect 14091 31298 14211 31336
rect 14091 31264 14114 31298
rect 14148 31264 14211 31298
rect 14091 31226 14211 31264
rect 14091 31192 14114 31226
rect 14148 31192 14211 31226
rect 14091 31154 14211 31192
rect 14091 31120 14114 31154
rect 14148 31120 14211 31154
rect 14091 31082 14211 31120
rect 14091 31048 14114 31082
rect 14148 31048 14211 31082
rect 14091 31010 14211 31048
rect 14091 30976 14114 31010
rect 14148 30976 14211 31010
rect 14091 30938 14211 30976
rect 14091 30904 14114 30938
rect 14148 30904 14211 30938
rect 14091 30866 14211 30904
rect 14091 30832 14114 30866
rect 14148 30832 14211 30866
rect 14091 30794 14211 30832
rect 14091 30760 14114 30794
rect 14148 30760 14211 30794
rect 14091 30722 14211 30760
rect 14091 30688 14114 30722
rect 14148 30688 14211 30722
rect 14091 30650 14211 30688
rect 14091 30616 14114 30650
rect 14148 30616 14211 30650
rect 14091 30578 14211 30616
rect 14091 30544 14114 30578
rect 14148 30544 14211 30578
rect 14091 30506 14211 30544
rect 14091 30472 14114 30506
rect 14148 30472 14211 30506
rect 14091 30434 14211 30472
rect 14091 30400 14114 30434
rect 14148 30400 14211 30434
rect 14091 30362 14211 30400
rect 14091 30328 14114 30362
rect 14148 30328 14211 30362
rect 14091 30290 14211 30328
rect 14091 30256 14114 30290
rect 14148 30256 14211 30290
rect 14091 30218 14211 30256
rect 14091 30184 14114 30218
rect 14148 30184 14211 30218
rect 14091 30146 14211 30184
rect 14091 30112 14114 30146
rect 14148 30112 14211 30146
rect 14091 30074 14211 30112
rect 14091 30040 14114 30074
rect 14148 30040 14211 30074
rect 14091 30002 14211 30040
rect 14091 29968 14114 30002
rect 14148 29968 14211 30002
rect 14091 29930 14211 29968
rect 14091 29896 14114 29930
rect 14148 29896 14211 29930
rect 14091 29858 14211 29896
rect 14091 29824 14114 29858
rect 14148 29824 14211 29858
rect 14091 29786 14211 29824
rect 14091 29752 14114 29786
rect 14148 29752 14211 29786
rect 14091 29714 14211 29752
rect 14091 29680 14114 29714
rect 14148 29680 14211 29714
rect 14091 29642 14211 29680
rect 14091 29608 14114 29642
rect 14148 29608 14211 29642
rect 14091 29570 14211 29608
rect 14091 29536 14114 29570
rect 14148 29536 14211 29570
rect 14091 29498 14211 29536
rect 14091 29464 14114 29498
rect 14148 29464 14211 29498
rect 14091 29426 14211 29464
rect 14091 29392 14114 29426
rect 14148 29392 14211 29426
rect 14091 29354 14211 29392
rect 14091 29320 14114 29354
rect 14148 29320 14211 29354
rect 14091 29282 14211 29320
rect 14091 29248 14114 29282
rect 14148 29248 14211 29282
rect 14091 29210 14211 29248
rect 14091 29176 14114 29210
rect 14148 29176 14211 29210
rect 14091 29138 14211 29176
rect 14091 29104 14114 29138
rect 14148 29104 14211 29138
rect 14091 29066 14211 29104
rect 14091 29032 14114 29066
rect 14148 29032 14211 29066
rect 14091 28994 14211 29032
rect 14091 28960 14114 28994
rect 14148 28960 14211 28994
rect 14091 28922 14211 28960
rect 14091 28888 14114 28922
rect 14148 28888 14211 28922
rect 14091 28850 14211 28888
rect 14091 28816 14114 28850
rect 14148 28816 14211 28850
rect 14091 28778 14211 28816
rect 14091 28744 14114 28778
rect 14148 28744 14211 28778
rect 14091 28706 14211 28744
rect 14091 28672 14114 28706
rect 14148 28672 14211 28706
rect 14091 28634 14211 28672
rect 14091 28600 14114 28634
rect 14148 28600 14211 28634
rect 14091 28562 14211 28600
rect 14091 28528 14114 28562
rect 14148 28528 14211 28562
rect 12915 28495 13556 28515
tri 2311 28289 2403 28381 se
rect 2403 28348 12596 28381
rect 2403 28289 4931 28348
rect 2311 28277 4931 28289
rect 7223 28277 7742 28348
rect 10034 28289 12596 28348
tri 12596 28289 12688 28381 sw
rect 10034 28277 12688 28289
rect 2311 28243 2443 28277
rect 2477 28243 2515 28277
rect 2549 28243 2587 28277
rect 2621 28243 2659 28277
rect 2693 28243 2731 28277
rect 2765 28243 2803 28277
rect 2837 28243 2875 28277
rect 2909 28243 2947 28277
rect 2981 28243 3019 28277
rect 3053 28243 3091 28277
rect 3125 28243 3163 28277
rect 3197 28243 3235 28277
rect 3269 28243 3307 28277
rect 3341 28243 3379 28277
rect 3413 28243 3451 28277
rect 3485 28243 3523 28277
rect 3557 28243 3595 28277
rect 3629 28243 3667 28277
rect 3701 28243 3739 28277
rect 3773 28243 3811 28277
rect 3845 28243 3883 28277
rect 3917 28243 3955 28277
rect 3989 28243 4027 28277
rect 4061 28243 4099 28277
rect 4133 28243 4171 28277
rect 4205 28243 4243 28277
rect 4277 28243 4315 28277
rect 4349 28243 4387 28277
rect 4421 28243 4459 28277
rect 4493 28243 4531 28277
rect 4565 28243 4603 28277
rect 4637 28243 4675 28277
rect 4709 28243 4747 28277
rect 4781 28243 4819 28277
rect 4853 28243 4891 28277
rect 4925 28243 4931 28277
rect 7229 28243 7267 28277
rect 7301 28243 7339 28277
rect 7373 28243 7411 28277
rect 7445 28243 7483 28277
rect 7517 28243 7555 28277
rect 7589 28243 7627 28277
rect 7661 28243 7699 28277
rect 7733 28243 7742 28277
rect 10037 28243 10075 28277
rect 10109 28243 10147 28277
rect 10181 28243 10219 28277
rect 10253 28243 10291 28277
rect 10325 28243 10363 28277
rect 10397 28243 10435 28277
rect 10469 28243 10507 28277
rect 10541 28243 10579 28277
rect 10613 28243 10651 28277
rect 10685 28243 10723 28277
rect 10757 28243 10795 28277
rect 10829 28243 10867 28277
rect 10901 28243 10939 28277
rect 10973 28243 11011 28277
rect 11045 28243 11083 28277
rect 11117 28243 11155 28277
rect 11189 28243 11227 28277
rect 11261 28243 11299 28277
rect 11333 28243 11371 28277
rect 11405 28243 11443 28277
rect 11477 28243 11515 28277
rect 11549 28243 11587 28277
rect 11621 28243 11659 28277
rect 11693 28243 11731 28277
rect 11765 28243 11803 28277
rect 11837 28243 11875 28277
rect 11909 28243 11947 28277
rect 11981 28243 12019 28277
rect 12053 28243 12091 28277
rect 12125 28243 12163 28277
rect 12197 28243 12235 28277
rect 12269 28243 12307 28277
rect 12341 28243 12379 28277
rect 12413 28243 12451 28277
rect 12485 28243 12523 28277
rect 12557 28243 12688 28277
rect 2311 28232 4931 28243
rect 7223 28232 7742 28243
rect 10034 28232 12688 28243
rect 2311 28203 12688 28232
rect 2311 28181 2479 28203
rect 2312 28169 2479 28181
rect 2513 28169 2551 28203
rect 2585 28169 2623 28203
rect 2657 28169 2695 28203
rect 2729 28169 2767 28203
rect 2801 28169 2839 28203
rect 2873 28169 2911 28203
rect 2945 28169 2983 28203
rect 3017 28169 3055 28203
rect 3089 28169 3127 28203
rect 3161 28169 3199 28203
rect 3233 28169 3271 28203
rect 3305 28169 3343 28203
rect 3377 28169 3415 28203
rect 3449 28169 3487 28203
rect 3521 28169 3559 28203
rect 3593 28169 3631 28203
rect 3665 28169 3703 28203
rect 3737 28169 3775 28203
rect 3809 28169 3847 28203
rect 3881 28169 3919 28203
rect 3953 28169 3991 28203
rect 4025 28169 4063 28203
rect 4097 28169 4135 28203
rect 4169 28169 4207 28203
rect 4241 28169 4279 28203
rect 4313 28169 4351 28203
rect 4385 28169 4423 28203
rect 4457 28169 4495 28203
rect 4529 28169 4567 28203
rect 4601 28169 4639 28203
rect 4673 28169 4711 28203
rect 4745 28169 4783 28203
rect 4817 28169 4855 28203
rect 4889 28169 4927 28203
rect 4961 28169 4999 28203
rect 5033 28169 5071 28203
rect 5105 28169 5143 28203
rect 5177 28169 5215 28203
rect 5249 28169 5287 28203
rect 5321 28169 5359 28203
rect 5393 28169 5431 28203
rect 5465 28169 5503 28203
rect 5537 28169 5575 28203
rect 5609 28169 5647 28203
rect 5681 28169 5719 28203
rect 5753 28169 5791 28203
rect 5825 28169 5863 28203
rect 5897 28169 5935 28203
rect 5969 28169 6007 28203
rect 6041 28169 6079 28203
rect 6113 28169 6151 28203
rect 6185 28169 6223 28203
rect 6257 28169 6295 28203
rect 6329 28169 6367 28203
rect 6401 28169 6439 28203
rect 6473 28169 6511 28203
rect 6545 28169 6583 28203
rect 6617 28169 6655 28203
rect 6689 28169 6727 28203
rect 6761 28169 6799 28203
rect 6833 28169 6871 28203
rect 6905 28169 6943 28203
rect 6977 28169 7015 28203
rect 7049 28169 7087 28203
rect 7121 28169 7159 28203
rect 7193 28169 7231 28203
rect 7265 28169 7303 28203
rect 7337 28169 7375 28203
rect 7409 28169 7447 28203
rect 7481 28169 7519 28203
rect 7553 28169 7591 28203
rect 7625 28169 7663 28203
rect 7697 28169 7735 28203
rect 7769 28169 7807 28203
rect 7841 28169 7879 28203
rect 7913 28169 7951 28203
rect 7985 28169 8023 28203
rect 8057 28169 8095 28203
rect 8129 28169 8167 28203
rect 8201 28169 8239 28203
rect 8273 28169 8311 28203
rect 8345 28169 8383 28203
rect 8417 28169 8455 28203
rect 8489 28169 8527 28203
rect 8561 28169 8599 28203
rect 8633 28169 8671 28203
rect 8705 28169 8743 28203
rect 8777 28169 8815 28203
rect 8849 28169 8887 28203
rect 8921 28169 8959 28203
rect 8993 28169 9031 28203
rect 9065 28169 9103 28203
rect 9137 28169 9175 28203
rect 9209 28169 9247 28203
rect 9281 28169 9319 28203
rect 9353 28169 9391 28203
rect 9425 28169 9463 28203
rect 9497 28169 9535 28203
rect 9569 28169 9607 28203
rect 9641 28169 9679 28203
rect 9713 28169 9751 28203
rect 9785 28169 9823 28203
rect 9857 28169 9895 28203
rect 9929 28169 9967 28203
rect 10001 28169 10039 28203
rect 10073 28169 10111 28203
rect 10145 28169 10183 28203
rect 10217 28169 10255 28203
rect 10289 28169 10327 28203
rect 10361 28169 10399 28203
rect 10433 28169 10471 28203
rect 10505 28169 10543 28203
rect 10577 28169 10615 28203
rect 10649 28169 10687 28203
rect 10721 28169 10759 28203
rect 10793 28169 10831 28203
rect 10865 28169 10903 28203
rect 10937 28169 10975 28203
rect 11009 28169 11047 28203
rect 11081 28169 11119 28203
rect 11153 28169 11191 28203
rect 11225 28169 11263 28203
rect 11297 28169 11335 28203
rect 11369 28169 11407 28203
rect 11441 28169 11479 28203
rect 11513 28169 11551 28203
rect 11585 28169 11623 28203
rect 11657 28169 11695 28203
rect 11729 28169 11767 28203
rect 11801 28169 11839 28203
rect 11873 28169 11911 28203
rect 11945 28169 11983 28203
rect 12017 28169 12055 28203
rect 12089 28169 12127 28203
rect 12161 28169 12199 28203
rect 12233 28169 12271 28203
rect 12305 28169 12343 28203
rect 12377 28169 12415 28203
rect 12449 28169 12487 28203
rect 12521 28169 12688 28203
rect 2312 28163 12688 28169
rect 2312 28104 2416 28163
tri 2416 28123 2456 28163 nw
tri 12544 28123 12584 28163 ne
rect 2312 28070 2376 28104
rect 2410 28070 2416 28104
rect 12584 28104 12688 28163
rect 2312 28032 2416 28070
rect 2312 27998 2376 28032
rect 2410 27998 2416 28032
rect 2312 27960 2416 27998
rect 2312 27926 2376 27960
rect 2410 27926 2416 27960
rect 2312 27888 2416 27926
rect 2312 27854 2376 27888
rect 2410 27854 2416 27888
tri 2480 28053 2500 28073 se
rect 2500 28053 12500 28073
tri 12500 28053 12520 28073 sw
rect 2480 28035 12520 28053
rect 2480 27919 2501 28035
rect 4473 28032 10492 28035
rect 12464 28032 12520 28035
rect 12485 27926 12520 28032
rect 4473 27919 10492 27926
rect 12464 27919 12520 27926
rect 2480 27905 12520 27919
tri 2480 27885 2500 27905 ne
rect 2500 27885 12500 27905
tri 12500 27885 12520 27905 nw
rect 12584 28070 12590 28104
rect 12624 28070 12688 28104
rect 12584 28032 12688 28070
rect 12584 27998 12590 28032
rect 12624 27998 12688 28032
rect 12584 27960 12688 27998
rect 12584 27926 12590 27960
rect 12624 27926 12688 27960
rect 12584 27888 12688 27926
rect 2312 27795 2416 27854
rect 12584 27854 12590 27888
rect 12624 27854 12688 27888
tri 2416 27795 2456 27835 sw
tri 12544 27795 12584 27835 se
rect 12584 27795 12688 27854
rect 2312 27789 12688 27795
rect 2312 27717 2479 27789
rect 2312 27683 2443 27717
rect 2477 27683 2479 27717
rect 12521 27717 12688 27789
rect 12521 27683 12523 27717
rect 12557 27683 12688 27717
rect 2312 27665 4931 27683
tri 2312 27565 2412 27665 ne
rect 2412 27616 4931 27665
rect 7223 27616 7742 27683
rect 10034 27665 12688 27683
rect 10034 27616 12588 27665
rect 2412 27565 12588 27616
tri 12588 27565 12688 27665 nw
rect 1651 27424 2085 27460
tri 2085 27424 2125 27464 sw
tri 12875 27424 12915 27464 se
rect 12915 27453 13023 28495
rect 13273 28296 13556 28495
tri 13556 28296 13775 28515 sw
rect 13273 27453 13775 28296
rect 12915 27424 13775 27453
rect 1651 27347 13775 27424
rect 1651 27230 1977 27347
tri 1651 27030 1851 27230 ne
rect 1851 27097 1977 27230
rect 13027 27230 13775 27347
rect 13027 27097 13149 27230
rect 1851 27030 13149 27097
tri 13149 27030 13349 27230 nw
rect 1111 26973 1153 27007
rect 1187 26973 1434 27007
rect 1111 26935 1434 26973
rect 1111 26901 1153 26935
rect 1187 26901 1434 26935
rect 1111 26863 1434 26901
rect 1111 26829 1153 26863
rect 1187 26829 1434 26863
rect 1111 26791 1434 26829
rect 1111 26757 1153 26791
rect 1187 26757 1434 26791
rect 1111 26719 1434 26757
rect 1111 26685 1153 26719
rect 1187 26685 1434 26719
rect 1111 26647 1434 26685
rect 1111 26613 1153 26647
rect 1187 26613 1434 26647
rect 1111 26575 1434 26613
rect 1111 26541 1153 26575
rect 1187 26541 1434 26575
rect 1111 26503 1434 26541
rect 1111 26469 1153 26503
rect 1187 26469 1434 26503
rect 1111 26431 1434 26469
rect 1111 26397 1153 26431
rect 1187 26397 1434 26431
rect 1111 26359 1434 26397
rect 1111 26325 1153 26359
rect 1187 26325 1434 26359
rect 1111 26287 1434 26325
rect 1111 26253 1153 26287
rect 1187 26253 1434 26287
rect 1111 26215 1434 26253
rect 1111 26181 1153 26215
rect 1187 26205 1434 26215
tri 1728 26205 2128 26605 se
rect 2128 26585 12848 26605
rect 2128 26205 2251 26585
rect 1187 26191 2251 26205
rect 12725 26205 12848 26585
tri 12848 26205 13248 26605 sw
rect 12725 26191 13248 26205
rect 1187 26181 13248 26191
rect 1111 26143 13248 26181
rect 1111 26109 1153 26143
rect 1187 26142 13248 26143
rect 1187 26109 2202 26142
rect 1111 26087 2202 26109
tri 2202 26102 2242 26142 nw
tri 12743 26102 12783 26142 ne
rect 1111 26071 1748 26087
rect 1111 26037 1153 26071
rect 1187 26037 1748 26071
rect 1111 25999 1748 26037
rect 1111 25965 1153 25999
rect 1187 25965 1748 25999
rect 1111 25927 1748 25965
rect 1111 25893 1153 25927
rect 1187 25893 1748 25927
rect 1111 25855 1748 25893
rect 1111 25821 1153 25855
rect 1187 25821 1748 25855
rect 1111 25783 1748 25821
rect 1111 25749 1153 25783
rect 1187 25749 1748 25783
rect 1111 25711 1748 25749
rect 1111 25677 1153 25711
rect 1187 25677 1748 25711
rect 1111 25639 1748 25677
rect 1111 25605 1153 25639
rect 1187 25605 1748 25639
rect 1111 25567 1748 25605
rect 1111 25533 1153 25567
rect 1187 25533 1748 25567
rect 1111 25495 1748 25533
rect 1111 25461 1153 25495
rect 1187 25461 1748 25495
rect 1111 25423 1748 25461
rect 1111 25389 1153 25423
rect 1187 25389 1748 25423
rect 1111 25351 1748 25389
rect 1111 25317 1153 25351
rect 1187 25333 1748 25351
rect 2142 25333 2202 26087
rect 12783 26087 13248 26142
tri 2383 26042 2406 26065 se
rect 2406 26042 12570 26065
tri 2320 25979 2383 26042 se
rect 2383 26038 12570 26042
rect 2383 25979 4925 26038
rect 2320 25922 4925 25979
rect 7217 25922 7749 26038
rect 10041 25979 12570 26038
tri 12570 25979 12656 26065 sw
rect 10041 25922 12656 25979
rect 2320 25909 12656 25922
rect 2320 25875 2503 25909
rect 2537 25875 2575 25909
rect 2609 25875 2647 25909
rect 2681 25875 2719 25909
rect 2753 25875 2791 25909
rect 2825 25875 2863 25909
rect 2897 25875 2935 25909
rect 2969 25875 3007 25909
rect 3041 25875 3079 25909
rect 3113 25875 3151 25909
rect 3185 25875 3223 25909
rect 3257 25875 3295 25909
rect 3329 25875 3367 25909
rect 3401 25875 3439 25909
rect 3473 25875 3511 25909
rect 3545 25875 3583 25909
rect 3617 25875 3655 25909
rect 3689 25875 3727 25909
rect 3761 25875 3799 25909
rect 3833 25875 3871 25909
rect 3905 25875 3943 25909
rect 3977 25875 4015 25909
rect 4049 25875 4087 25909
rect 4121 25875 4159 25909
rect 4193 25875 4231 25909
rect 4265 25875 4303 25909
rect 4337 25875 4375 25909
rect 4409 25875 4447 25909
rect 4481 25875 4519 25909
rect 4553 25875 4591 25909
rect 4625 25875 4663 25909
rect 4697 25875 4735 25909
rect 4769 25875 4807 25909
rect 4841 25875 4879 25909
rect 4913 25875 4951 25909
rect 4985 25875 5023 25909
rect 5057 25875 5095 25909
rect 5129 25875 5167 25909
rect 5201 25875 5239 25909
rect 5273 25875 5311 25909
rect 5345 25875 5383 25909
rect 5417 25875 5455 25909
rect 5489 25875 5527 25909
rect 5561 25875 5599 25909
rect 5633 25875 5671 25909
rect 5705 25875 5743 25909
rect 5777 25875 5815 25909
rect 5849 25875 5887 25909
rect 5921 25875 5959 25909
rect 5993 25875 6031 25909
rect 6065 25875 6103 25909
rect 6137 25875 6175 25909
rect 6209 25875 6247 25909
rect 6281 25875 6319 25909
rect 6353 25875 6391 25909
rect 6425 25875 6463 25909
rect 6497 25875 6535 25909
rect 6569 25875 6607 25909
rect 6641 25875 6679 25909
rect 6713 25875 6751 25909
rect 6785 25875 6823 25909
rect 6857 25875 6895 25909
rect 6929 25875 6967 25909
rect 7001 25875 7039 25909
rect 7073 25875 7111 25909
rect 7145 25875 7183 25909
rect 7217 25875 7255 25909
rect 7289 25875 7327 25909
rect 7361 25875 7399 25909
rect 7433 25875 7471 25909
rect 7505 25875 7543 25909
rect 7577 25875 7615 25909
rect 7649 25875 7687 25909
rect 7721 25875 7759 25909
rect 7793 25875 7831 25909
rect 7865 25875 7903 25909
rect 7937 25875 7975 25909
rect 8009 25875 8047 25909
rect 8081 25875 8119 25909
rect 8153 25875 8191 25909
rect 8225 25875 8263 25909
rect 8297 25875 8335 25909
rect 8369 25875 8407 25909
rect 8441 25875 8479 25909
rect 8513 25875 8551 25909
rect 8585 25875 8623 25909
rect 8657 25875 8695 25909
rect 8729 25875 8767 25909
rect 8801 25875 8839 25909
rect 8873 25875 8911 25909
rect 8945 25875 8983 25909
rect 9017 25875 9055 25909
rect 9089 25875 9127 25909
rect 9161 25875 9199 25909
rect 9233 25875 9271 25909
rect 9305 25875 9343 25909
rect 9377 25875 9415 25909
rect 9449 25875 9487 25909
rect 9521 25875 9559 25909
rect 9593 25875 9631 25909
rect 9665 25875 9703 25909
rect 9737 25875 9775 25909
rect 9809 25875 9847 25909
rect 9881 25875 9919 25909
rect 9953 25875 9991 25909
rect 10025 25875 10063 25909
rect 10097 25875 10135 25909
rect 10169 25875 10207 25909
rect 10241 25875 10279 25909
rect 10313 25875 10351 25909
rect 10385 25875 10423 25909
rect 10457 25875 10495 25909
rect 10529 25875 10567 25909
rect 10601 25875 10639 25909
rect 10673 25875 10711 25909
rect 10745 25875 10783 25909
rect 10817 25875 10855 25909
rect 10889 25875 10927 25909
rect 10961 25875 10999 25909
rect 11033 25875 11071 25909
rect 11105 25875 11143 25909
rect 11177 25875 11215 25909
rect 11249 25875 11287 25909
rect 11321 25875 11359 25909
rect 11393 25875 11431 25909
rect 11465 25875 11503 25909
rect 11537 25875 11575 25909
rect 11609 25875 11647 25909
rect 11681 25875 11719 25909
rect 11753 25875 11791 25909
rect 11825 25875 11863 25909
rect 11897 25875 11935 25909
rect 11969 25875 12007 25909
rect 12041 25875 12079 25909
rect 12113 25875 12151 25909
rect 12185 25875 12223 25909
rect 12257 25875 12295 25909
rect 12329 25875 12367 25909
rect 12401 25875 12439 25909
rect 12473 25875 12656 25909
rect 2320 25869 12656 25875
rect 2320 25796 2426 25869
tri 2426 25829 2466 25869 nw
tri 12510 25829 12550 25869 ne
rect 2320 25762 2386 25796
rect 2420 25762 2426 25796
rect 2320 25724 2426 25762
rect 2320 25690 2386 25724
rect 2420 25690 2426 25724
rect 2320 25652 2426 25690
rect 2320 25618 2386 25652
rect 2420 25618 2426 25652
rect 2320 25545 2426 25618
tri 2468 25781 2488 25801 se
rect 2488 25781 12488 25801
tri 12488 25781 12508 25801 sw
rect 2468 25772 12508 25781
rect 2468 25760 2538 25772
rect 4446 25760 10520 25772
rect 12428 25760 12508 25772
rect 2468 25654 2503 25760
rect 12473 25654 12508 25760
rect 2468 25633 12508 25654
tri 2468 25613 2488 25633 ne
rect 2488 25613 12488 25633
tri 12488 25613 12508 25633 nw
rect 12550 25796 12656 25869
rect 12550 25762 12556 25796
rect 12590 25762 12656 25796
rect 12550 25724 12656 25762
rect 12550 25690 12556 25724
rect 12590 25690 12656 25724
rect 12550 25652 12656 25690
rect 12550 25618 12556 25652
rect 12590 25618 12656 25652
tri 2426 25545 2466 25585 sw
tri 12510 25545 12550 25585 se
rect 12550 25545 12656 25618
rect 2320 25539 12656 25545
rect 2320 25533 2503 25539
rect 2318 25505 2503 25533
rect 2537 25505 2575 25539
rect 2609 25505 2647 25539
rect 2681 25505 2719 25539
rect 2753 25505 2791 25539
rect 2825 25505 2863 25539
rect 2897 25505 2935 25539
rect 2969 25505 3007 25539
rect 3041 25505 3079 25539
rect 3113 25505 3151 25539
rect 3185 25505 3223 25539
rect 3257 25505 3295 25539
rect 3329 25505 3367 25539
rect 3401 25505 3439 25539
rect 3473 25505 3511 25539
rect 3545 25505 3583 25539
rect 3617 25505 3655 25539
rect 3689 25505 3727 25539
rect 3761 25505 3799 25539
rect 3833 25505 3871 25539
rect 3905 25505 3943 25539
rect 3977 25505 4015 25539
rect 4049 25505 4087 25539
rect 4121 25505 4159 25539
rect 4193 25505 4231 25539
rect 4265 25505 4303 25539
rect 4337 25505 4375 25539
rect 4409 25505 4447 25539
rect 4481 25505 4519 25539
rect 4553 25505 4591 25539
rect 4625 25505 4663 25539
rect 4697 25505 4735 25539
rect 4769 25505 4807 25539
rect 4841 25505 4879 25539
rect 4913 25506 4951 25539
rect 4985 25506 5023 25539
rect 5057 25506 5095 25539
rect 5129 25506 5167 25539
rect 5201 25506 5239 25539
rect 5273 25506 5311 25539
rect 5345 25506 5383 25539
rect 5417 25506 5455 25539
rect 5489 25506 5527 25539
rect 5561 25506 5599 25539
rect 5633 25506 5671 25539
rect 5705 25506 5743 25539
rect 5777 25506 5815 25539
rect 5849 25506 5887 25539
rect 5921 25506 5959 25539
rect 5993 25506 6031 25539
rect 6065 25506 6103 25539
rect 6137 25506 6175 25539
rect 6209 25506 6247 25539
rect 6281 25506 6319 25539
rect 6353 25506 6391 25539
rect 6425 25506 6463 25539
rect 6497 25506 6535 25539
rect 6569 25506 6607 25539
rect 6641 25506 6679 25539
rect 6713 25506 6751 25539
rect 6785 25506 6823 25539
rect 6857 25506 6895 25539
rect 6929 25506 6967 25539
rect 7001 25506 7039 25539
rect 7073 25506 7111 25539
rect 7145 25506 7183 25539
rect 4913 25505 4925 25506
rect 7217 25505 7255 25539
rect 7289 25505 7327 25539
rect 7361 25505 7399 25539
rect 7433 25505 7471 25539
rect 7505 25505 7543 25539
rect 7577 25505 7615 25539
rect 7649 25505 7687 25539
rect 7721 25506 7759 25539
rect 7793 25506 7831 25539
rect 7865 25506 7903 25539
rect 7937 25506 7975 25539
rect 8009 25506 8047 25539
rect 8081 25506 8119 25539
rect 8153 25506 8191 25539
rect 8225 25506 8263 25539
rect 8297 25506 8335 25539
rect 8369 25506 8407 25539
rect 8441 25506 8479 25539
rect 8513 25506 8551 25539
rect 8585 25506 8623 25539
rect 8657 25506 8695 25539
rect 8729 25506 8767 25539
rect 8801 25506 8839 25539
rect 8873 25506 8911 25539
rect 8945 25506 8983 25539
rect 9017 25506 9055 25539
rect 9089 25506 9127 25539
rect 9161 25506 9199 25539
rect 9233 25506 9271 25539
rect 9305 25506 9343 25539
rect 9377 25506 9415 25539
rect 9449 25506 9487 25539
rect 9521 25506 9559 25539
rect 9593 25506 9631 25539
rect 9665 25506 9703 25539
rect 9737 25506 9775 25539
rect 9809 25506 9847 25539
rect 9881 25506 9919 25539
rect 9953 25506 9991 25539
rect 10025 25506 10063 25539
rect 7721 25505 7749 25506
rect 10041 25505 10063 25506
rect 10097 25505 10135 25539
rect 10169 25505 10207 25539
rect 10241 25505 10279 25539
rect 10313 25505 10351 25539
rect 10385 25505 10423 25539
rect 10457 25505 10495 25539
rect 10529 25505 10567 25539
rect 10601 25505 10639 25539
rect 10673 25505 10711 25539
rect 10745 25505 10783 25539
rect 10817 25505 10855 25539
rect 10889 25505 10927 25539
rect 10961 25505 10999 25539
rect 11033 25505 11071 25539
rect 11105 25505 11143 25539
rect 11177 25505 11215 25539
rect 11249 25505 11287 25539
rect 11321 25505 11359 25539
rect 11393 25505 11431 25539
rect 11465 25505 11503 25539
rect 11537 25505 11575 25539
rect 11609 25505 11647 25539
rect 11681 25505 11719 25539
rect 11753 25505 11791 25539
rect 11825 25505 11863 25539
rect 11897 25505 11935 25539
rect 11969 25505 12007 25539
rect 12041 25505 12079 25539
rect 12113 25505 12151 25539
rect 12185 25505 12223 25539
rect 12257 25505 12295 25539
rect 12329 25505 12367 25539
rect 12401 25505 12439 25539
rect 12473 25505 12656 25539
rect 2318 25441 4925 25505
tri 2318 25361 2398 25441 ne
rect 2398 25390 4925 25441
rect 7217 25390 7749 25505
rect 10041 25441 12656 25505
rect 10041 25390 12574 25441
rect 2398 25361 12574 25390
tri 12574 25361 12654 25441 nw
rect 1187 25317 2202 25333
rect 12783 25333 12834 26087
rect 13228 25333 13248 26087
rect 1111 25283 2202 25317
tri 2202 25283 2242 25323 sw
tri 12743 25283 12783 25323 se
rect 12783 25283 13248 25333
rect 1111 25279 13248 25283
rect 1111 25245 1153 25279
rect 1187 25245 13248 25279
rect 1111 25229 13248 25245
rect 1111 25215 2251 25229
rect 1111 25207 1229 25215
rect 1111 25173 1153 25207
rect 1187 25173 1229 25207
rect 1111 25135 1229 25173
rect 1111 25101 1153 25135
rect 1187 25101 1229 25135
rect 1111 25063 1229 25101
rect 1111 25029 1153 25063
rect 1187 25029 1229 25063
rect 1111 24991 1229 25029
rect 1111 24957 1153 24991
rect 1187 24957 1229 24991
rect 1111 24919 1229 24957
rect 1111 24885 1153 24919
rect 1187 24885 1229 24919
rect 1111 24847 1229 24885
rect 1111 24813 1153 24847
rect 1187 24813 1229 24847
tri 1728 24815 2128 25215 ne
rect 2128 24835 2251 25215
rect 12725 25215 13248 25229
rect 12725 24835 12848 25215
rect 2128 24815 12848 24835
tri 12848 24815 13248 25215 nw
rect 1111 24775 1229 24813
rect 1111 24741 1153 24775
rect 1187 24741 1229 24775
rect 1111 24703 1229 24741
rect 1111 24669 1153 24703
rect 1187 24669 1229 24703
rect 1111 24631 1229 24669
rect 1111 24597 1153 24631
rect 1187 24597 1229 24631
rect 1111 24559 1229 24597
rect 1111 24525 1153 24559
rect 1187 24525 1229 24559
rect 13519 24556 13775 27230
tri 4857 24530 4883 24556 se
rect 4883 24530 13775 24556
rect 1111 24487 1229 24525
rect 1111 24453 1153 24487
rect 1187 24453 1229 24487
rect 1111 24415 1229 24453
rect 1111 24381 1153 24415
rect 1187 24381 1229 24415
rect 1111 24343 1229 24381
rect 1111 24309 1153 24343
rect 1187 24309 1229 24343
rect 1111 24271 1229 24309
rect 1111 24237 1153 24271
rect 1187 24237 1229 24271
rect 1111 24199 1229 24237
rect 1111 24165 1153 24199
rect 1187 24165 1229 24199
rect 1111 24127 1229 24165
rect 1111 24093 1153 24127
rect 1187 24093 1229 24127
rect 1111 24055 1229 24093
rect 1111 24021 1153 24055
rect 1187 24021 1229 24055
rect 1111 23983 1229 24021
rect 1111 23949 1153 23983
rect 1187 23949 1229 23983
rect 1111 23911 1229 23949
rect 1111 23877 1153 23911
rect 1187 23877 1229 23911
rect 1111 23839 1229 23877
rect 1111 23805 1153 23839
rect 1187 23805 1229 23839
rect 1111 23767 1229 23805
rect 1111 23733 1153 23767
rect 1187 23733 1229 23767
rect 1111 23695 1229 23733
rect 1111 23661 1153 23695
rect 1187 23661 1229 23695
rect 1111 23623 1229 23661
tri 4683 24356 4857 24530 se
rect 4857 24502 13775 24530
rect 4857 24356 4937 24502
rect 4683 23828 4937 24356
tri 4683 23628 4883 23828 ne
rect 4883 23682 4937 23828
rect 7229 23682 7736 24502
rect 10028 24054 13775 24502
rect 10028 23682 13349 24054
rect 4883 23628 13349 23682
tri 13349 23628 13775 24054 nw
rect 14091 28490 14211 28528
rect 14091 28456 14114 28490
rect 14148 28456 14211 28490
rect 14091 28418 14211 28456
rect 14091 28384 14114 28418
rect 14148 28384 14211 28418
rect 14091 28346 14211 28384
rect 14091 28312 14114 28346
rect 14148 28312 14211 28346
rect 14091 28274 14211 28312
rect 14091 28240 14114 28274
rect 14148 28240 14211 28274
rect 14091 28202 14211 28240
rect 14091 28168 14114 28202
rect 14148 28168 14211 28202
rect 14091 28130 14211 28168
rect 14091 28096 14114 28130
rect 14148 28096 14211 28130
rect 14091 28058 14211 28096
rect 14091 28024 14114 28058
rect 14148 28024 14211 28058
rect 14091 27986 14211 28024
rect 14091 27952 14114 27986
rect 14148 27952 14211 27986
rect 14091 27914 14211 27952
rect 14091 27880 14114 27914
rect 14148 27880 14211 27914
rect 14091 27842 14211 27880
rect 14091 27808 14114 27842
rect 14148 27808 14211 27842
rect 14091 27770 14211 27808
rect 14091 27736 14114 27770
rect 14148 27736 14211 27770
rect 14091 27698 14211 27736
rect 14091 27664 14114 27698
rect 14148 27664 14211 27698
rect 14091 27626 14211 27664
rect 14091 27592 14114 27626
rect 14148 27592 14211 27626
rect 14091 27554 14211 27592
rect 14091 27520 14114 27554
rect 14148 27520 14211 27554
rect 14091 27482 14211 27520
rect 14091 27448 14114 27482
rect 14148 27448 14211 27482
rect 14091 27410 14211 27448
rect 14091 27376 14114 27410
rect 14148 27376 14211 27410
rect 14091 27338 14211 27376
rect 14091 27304 14114 27338
rect 14148 27304 14211 27338
rect 14091 27266 14211 27304
rect 14091 27232 14114 27266
rect 14148 27232 14211 27266
rect 14091 27194 14211 27232
rect 14091 27160 14114 27194
rect 14148 27160 14211 27194
rect 14091 27122 14211 27160
rect 14091 27088 14114 27122
rect 14148 27088 14211 27122
rect 14091 27050 14211 27088
rect 14091 27016 14114 27050
rect 14148 27016 14211 27050
rect 14091 26978 14211 27016
rect 14091 26944 14114 26978
rect 14148 26944 14211 26978
rect 14091 26906 14211 26944
rect 14091 26872 14114 26906
rect 14148 26872 14211 26906
rect 14091 26834 14211 26872
rect 14091 26800 14114 26834
rect 14148 26800 14211 26834
rect 14091 26762 14211 26800
rect 14091 26728 14114 26762
rect 14148 26728 14211 26762
rect 14091 26690 14211 26728
rect 14091 26656 14114 26690
rect 14148 26656 14211 26690
rect 14091 26618 14211 26656
rect 14091 26584 14114 26618
rect 14148 26584 14211 26618
rect 14091 26546 14211 26584
rect 14091 26512 14114 26546
rect 14148 26512 14211 26546
rect 14091 26474 14211 26512
rect 14091 26440 14114 26474
rect 14148 26440 14211 26474
rect 14091 26402 14211 26440
rect 14091 26368 14114 26402
rect 14148 26368 14211 26402
rect 14091 26330 14211 26368
rect 14091 26296 14114 26330
rect 14148 26296 14211 26330
rect 14091 26258 14211 26296
rect 14091 26224 14114 26258
rect 14148 26224 14211 26258
rect 14091 26186 14211 26224
rect 14091 26152 14114 26186
rect 14148 26152 14211 26186
rect 14091 26114 14211 26152
rect 14091 26080 14114 26114
rect 14148 26080 14211 26114
rect 14091 26042 14211 26080
rect 14091 26008 14114 26042
rect 14148 26008 14211 26042
rect 14091 25970 14211 26008
rect 14091 25936 14114 25970
rect 14148 25936 14211 25970
rect 14091 25898 14211 25936
rect 14091 25864 14114 25898
rect 14148 25864 14211 25898
rect 14091 25826 14211 25864
rect 14091 25792 14114 25826
rect 14148 25792 14211 25826
rect 14091 25754 14211 25792
rect 14091 25720 14114 25754
rect 14148 25720 14211 25754
rect 14091 25682 14211 25720
rect 14091 25648 14114 25682
rect 14148 25648 14211 25682
rect 14091 25610 14211 25648
rect 14091 25576 14114 25610
rect 14148 25576 14211 25610
rect 14091 25538 14211 25576
rect 14091 25504 14114 25538
rect 14148 25504 14211 25538
rect 14091 25466 14211 25504
rect 14091 25432 14114 25466
rect 14148 25432 14211 25466
rect 14091 25394 14211 25432
rect 14091 25360 14114 25394
rect 14148 25360 14211 25394
rect 14091 25322 14211 25360
rect 14091 25288 14114 25322
rect 14148 25288 14211 25322
rect 14091 25250 14211 25288
rect 14091 25216 14114 25250
rect 14148 25216 14211 25250
rect 14091 25178 14211 25216
rect 14091 25144 14114 25178
rect 14148 25144 14211 25178
rect 14091 25106 14211 25144
rect 14091 25072 14114 25106
rect 14148 25072 14211 25106
rect 14091 25034 14211 25072
rect 14091 25000 14114 25034
rect 14148 25000 14211 25034
rect 14091 24962 14211 25000
rect 14091 24928 14114 24962
rect 14148 24928 14211 24962
rect 14091 24890 14211 24928
rect 14091 24856 14114 24890
rect 14148 24856 14211 24890
rect 14091 24818 14211 24856
rect 14091 24784 14114 24818
rect 14148 24784 14211 24818
rect 14091 24746 14211 24784
rect 14091 24712 14114 24746
rect 14148 24712 14211 24746
rect 14091 24674 14211 24712
rect 14091 24640 14114 24674
rect 14148 24640 14211 24674
rect 14091 24602 14211 24640
rect 14091 24568 14114 24602
rect 14148 24568 14211 24602
rect 14091 24530 14211 24568
rect 14091 24496 14114 24530
rect 14148 24496 14211 24530
rect 14091 24458 14211 24496
rect 14091 24424 14114 24458
rect 14148 24424 14211 24458
rect 14091 24386 14211 24424
rect 14091 24352 14114 24386
rect 14148 24352 14211 24386
rect 14091 24314 14211 24352
rect 14091 24280 14114 24314
rect 14148 24280 14211 24314
rect 14091 24242 14211 24280
rect 14091 24208 14114 24242
rect 14148 24208 14211 24242
rect 14091 24170 14211 24208
rect 14091 24136 14114 24170
rect 14148 24136 14211 24170
rect 14091 24098 14211 24136
rect 14091 24064 14114 24098
rect 14148 24064 14211 24098
rect 14091 24026 14211 24064
rect 14091 23992 14114 24026
rect 14148 23992 14211 24026
rect 14091 23954 14211 23992
rect 14091 23920 14114 23954
rect 14148 23920 14211 23954
rect 14091 23882 14211 23920
rect 14091 23848 14114 23882
rect 14148 23848 14211 23882
rect 14091 23810 14211 23848
rect 14091 23776 14114 23810
rect 14148 23776 14211 23810
rect 14091 23738 14211 23776
rect 14091 23704 14114 23738
rect 14148 23704 14211 23738
rect 14091 23666 14211 23704
rect 14091 23632 14114 23666
rect 14148 23632 14211 23666
rect 1111 23589 1153 23623
rect 1187 23589 1229 23623
rect 1111 23551 1229 23589
rect 1111 23517 1153 23551
rect 1187 23517 1229 23551
rect 1111 23479 1229 23517
rect 1111 23445 1153 23479
rect 1187 23445 1229 23479
rect 1111 23407 1229 23445
rect 14091 23594 14211 23632
rect 14091 23560 14114 23594
rect 14148 23560 14211 23594
rect 14091 23522 14211 23560
rect 14091 23488 14114 23522
rect 14148 23488 14211 23522
rect 14091 23450 14211 23488
rect 1111 23373 1153 23407
rect 1187 23373 1229 23407
rect 1111 23335 1229 23373
rect 1111 23301 1153 23335
rect 1187 23301 1229 23335
rect 1111 23263 1229 23301
rect 1111 23229 1153 23263
rect 1187 23229 1229 23263
rect 1111 23191 1229 23229
rect 1111 23157 1153 23191
rect 1187 23157 1229 23191
rect 1111 23119 1229 23157
rect 1111 23085 1153 23119
rect 1187 23085 1229 23119
rect 1111 23047 1229 23085
rect 1111 23013 1153 23047
rect 1187 23013 1229 23047
rect 1111 22975 1229 23013
rect 1111 22941 1153 22975
rect 1187 22941 1229 22975
rect 1111 22903 1229 22941
rect 1111 22869 1153 22903
rect 1187 22869 1229 22903
rect 1111 22831 1229 22869
rect 1111 22797 1153 22831
rect 1187 22797 1229 22831
rect 1111 22759 1229 22797
rect 1111 22725 1153 22759
rect 1187 22725 1229 22759
rect 1111 22687 1229 22725
rect 1111 22653 1153 22687
rect 1187 22653 1229 22687
rect 1111 22615 1229 22653
rect 1111 22581 1153 22615
rect 1187 22581 1229 22615
rect 1111 22543 1229 22581
rect 1111 22509 1153 22543
rect 1187 22509 1229 22543
rect 1111 22471 1229 22509
rect 1111 22437 1153 22471
rect 1187 22437 1229 22471
rect 1111 22399 1229 22437
rect 1111 22365 1153 22399
rect 1187 22365 1229 22399
rect 1111 22327 1229 22365
rect 1111 22293 1153 22327
rect 1187 22293 1229 22327
rect 1111 22255 1229 22293
rect 1111 22221 1153 22255
rect 1187 22221 1229 22255
rect 1111 22183 1229 22221
rect 1111 22149 1153 22183
rect 1187 22149 1229 22183
rect 1111 22111 1229 22149
rect 1111 22077 1153 22111
rect 1187 22077 1229 22111
rect 1111 22039 1229 22077
rect 1111 22005 1153 22039
rect 1187 22005 1229 22039
rect 1111 21967 1229 22005
rect 1111 21933 1153 21967
rect 1187 21933 1229 21967
rect 1111 21895 1229 21933
rect 1111 21861 1153 21895
rect 1187 21861 1229 21895
rect 1111 21823 1229 21861
rect 1111 21789 1153 21823
rect 1187 21789 1229 21823
rect 1111 21751 1229 21789
rect 1111 21717 1153 21751
rect 1187 21717 1229 21751
rect 1111 21679 1229 21717
rect 1111 21645 1153 21679
rect 1187 21645 1229 21679
rect 1111 21607 1229 21645
rect 1111 21573 1153 21607
rect 1187 21573 1229 21607
rect 1111 21535 1229 21573
rect 1111 21501 1153 21535
rect 1187 21501 1229 21535
rect 1111 21463 1229 21501
rect 1111 21429 1153 21463
rect 1187 21429 1229 21463
rect 1111 21391 1229 21429
rect 1111 21357 1153 21391
rect 1187 21357 1229 21391
rect 1111 21319 1229 21357
rect 1111 21285 1153 21319
rect 1187 21285 1229 21319
rect 1111 21247 1229 21285
rect 1111 21213 1153 21247
rect 1187 21213 1229 21247
rect 1111 21175 1229 21213
rect 1111 21141 1153 21175
rect 1187 21141 1229 21175
rect 1111 21103 1229 21141
rect 1111 21069 1153 21103
rect 1187 21069 1229 21103
rect 1111 21031 1229 21069
rect 1111 20997 1153 21031
rect 1187 20997 1229 21031
rect 1111 20959 1229 20997
rect 1111 20925 1153 20959
rect 1187 20925 1229 20959
rect 1111 20887 1229 20925
rect 1111 20853 1153 20887
rect 1187 20853 1229 20887
rect 1111 20815 1229 20853
rect 1111 20781 1153 20815
rect 1187 20781 1229 20815
rect 1111 20743 1229 20781
rect 1111 20709 1153 20743
rect 1187 20709 1229 20743
rect 1111 20671 1229 20709
rect 1111 20637 1153 20671
rect 1187 20637 1229 20671
rect 1111 20599 1229 20637
rect 1111 20565 1153 20599
rect 1187 20565 1229 20599
rect 1111 20527 1229 20565
rect 1111 20493 1153 20527
rect 1187 20493 1229 20527
rect 1111 20455 1229 20493
rect 1111 20421 1153 20455
rect 1187 20421 1229 20455
rect 1111 20383 1229 20421
rect 1111 20349 1153 20383
rect 1187 20349 1229 20383
rect 1111 20311 1229 20349
rect 1111 20277 1153 20311
rect 1187 20277 1229 20311
rect 1111 20239 1229 20277
rect 1111 20205 1153 20239
rect 1187 20205 1229 20239
rect 1111 20167 1229 20205
rect 1111 20133 1153 20167
rect 1187 20133 1229 20167
rect 1111 20095 1229 20133
rect 1111 20061 1153 20095
rect 1187 20061 1229 20095
rect 1111 20023 1229 20061
rect 1111 19989 1153 20023
rect 1187 19989 1229 20023
rect 1111 19951 1229 19989
rect 1111 19917 1153 19951
rect 1187 19917 1229 19951
rect 1111 19879 1229 19917
rect 1111 19845 1153 19879
rect 1187 19845 1229 19879
rect 1111 19807 1229 19845
rect 1111 19773 1153 19807
rect 1187 19773 1229 19807
rect 1111 19735 1229 19773
rect 1111 19701 1153 19735
rect 1187 19701 1229 19735
rect 1111 19663 1229 19701
rect 1111 19629 1153 19663
rect 1187 19629 1229 19663
rect 1111 19591 1229 19629
rect 1111 19557 1153 19591
rect 1187 19557 1229 19591
rect 1111 19519 1229 19557
rect 1111 19485 1153 19519
rect 1187 19485 1229 19519
rect 1111 19447 1229 19485
rect 1111 19413 1153 19447
rect 1187 19413 1229 19447
rect 1111 19375 1229 19413
rect 1111 19341 1153 19375
rect 1187 19341 1229 19375
rect 1111 19303 1229 19341
rect 1111 19269 1153 19303
rect 1187 19269 1229 19303
rect 1111 19231 1229 19269
rect 1111 19197 1153 19231
rect 1187 19197 1229 19231
rect 1111 19159 1229 19197
rect 1111 19125 1153 19159
rect 1187 19125 1229 19159
rect 1111 19087 1229 19125
rect 1111 19053 1153 19087
rect 1187 19053 1229 19087
rect 1111 19015 1229 19053
rect 1111 18981 1153 19015
rect 1187 18981 1229 19015
rect 1111 18943 1229 18981
rect 1111 18909 1153 18943
rect 1187 18909 1229 18943
rect 1111 18871 1229 18909
rect 1111 18837 1153 18871
rect 1187 18837 1229 18871
rect 1111 18799 1229 18837
rect 1111 18765 1153 18799
rect 1187 18765 1229 18799
rect 1111 18727 1229 18765
rect 1111 18693 1153 18727
rect 1187 18693 1229 18727
rect 1111 18655 1229 18693
rect 1111 18621 1153 18655
rect 1187 18621 1229 18655
rect 1111 18583 1229 18621
rect 1111 18549 1153 18583
rect 1187 18549 1229 18583
rect 1111 18511 1229 18549
rect 1111 18477 1153 18511
rect 1187 18477 1229 18511
rect 1111 18439 1229 18477
rect 1111 18405 1153 18439
rect 1187 18405 1229 18439
rect 1111 18367 1229 18405
rect 1111 18333 1153 18367
rect 1187 18333 1229 18367
rect 1111 18295 1229 18333
rect 1111 18261 1153 18295
rect 1187 18261 1229 18295
rect 1111 18223 1229 18261
rect 1111 18189 1153 18223
rect 1187 18189 1229 18223
rect 1111 18151 1229 18189
rect 1111 18117 1153 18151
rect 1187 18117 1229 18151
rect 1111 18079 1229 18117
rect 1111 18045 1153 18079
rect 1187 18045 1229 18079
rect 1111 18007 1229 18045
rect 1111 17973 1153 18007
rect 1187 17973 1229 18007
rect 1111 17935 1229 17973
rect 1111 17901 1153 17935
rect 1187 17901 1229 17935
rect 1111 17863 1229 17901
rect 1111 17829 1153 17863
rect 1187 17829 1229 17863
rect 1111 17791 1229 17829
rect 1111 17757 1153 17791
rect 1187 17757 1229 17791
rect 1111 17719 1229 17757
rect 1111 17685 1153 17719
rect 1187 17685 1229 17719
rect 1111 17647 1229 17685
rect 1111 17613 1153 17647
rect 1187 17613 1229 17647
rect 1111 17575 1229 17613
rect 1111 17541 1153 17575
rect 1187 17541 1229 17575
rect 1111 17503 1229 17541
rect 1111 17469 1153 17503
rect 1187 17469 1229 17503
rect 1111 17431 1229 17469
rect 1111 17397 1153 17431
rect 1187 17397 1229 17431
rect 1111 17359 1229 17397
rect 1111 17325 1153 17359
rect 1187 17325 1229 17359
rect 1111 17287 1229 17325
rect 1111 17253 1153 17287
rect 1187 17253 1229 17287
rect 1111 17215 1229 17253
rect 1111 17181 1153 17215
rect 1187 17181 1229 17215
rect 1111 17143 1229 17181
rect 1111 17109 1153 17143
rect 1187 17109 1229 17143
rect 1111 17071 1229 17109
rect 1111 17037 1153 17071
rect 1187 17037 1229 17071
rect 1111 16999 1229 17037
rect 1111 16965 1153 16999
rect 1187 16965 1229 16999
rect 1111 16927 1229 16965
rect 1111 16893 1153 16927
rect 1187 16893 1229 16927
rect 1111 16855 1229 16893
rect 1111 16821 1153 16855
rect 1187 16821 1229 16855
rect 1111 16783 1229 16821
rect 1111 16749 1153 16783
rect 1187 16749 1229 16783
rect 1111 16711 1229 16749
rect 1111 16677 1153 16711
rect 1187 16677 1229 16711
rect 1111 16639 1229 16677
rect 1111 16605 1153 16639
rect 1187 16605 1229 16639
rect 1111 16567 1229 16605
rect 1111 16533 1153 16567
rect 1187 16533 1229 16567
rect 1111 16495 1229 16533
rect 1111 16461 1153 16495
rect 1187 16461 1229 16495
rect 1111 16423 1229 16461
rect 1111 16389 1153 16423
rect 1187 16389 1229 16423
rect 1111 16351 1229 16389
rect 1111 16317 1153 16351
rect 1187 16317 1229 16351
rect 1111 16279 1229 16317
rect 1111 16245 1153 16279
rect 1187 16245 1229 16279
rect 1111 16207 1229 16245
rect 1111 16173 1153 16207
rect 1187 16173 1229 16207
rect 1111 16135 1229 16173
rect 1111 16101 1153 16135
rect 1187 16101 1229 16135
rect 1111 16063 1229 16101
rect 1111 16029 1153 16063
rect 1187 16029 1229 16063
rect 1111 15991 1229 16029
rect 1111 15957 1153 15991
rect 1187 15957 1229 15991
rect 1111 15919 1229 15957
rect 1111 15885 1153 15919
rect 1187 15885 1229 15919
rect 1111 15847 1229 15885
rect 1111 15813 1153 15847
rect 1187 15813 1229 15847
rect 1111 15775 1229 15813
rect 1111 15741 1153 15775
rect 1187 15741 1229 15775
rect 1111 15703 1229 15741
rect 1111 15669 1153 15703
rect 1187 15669 1229 15703
rect 1111 15631 1229 15669
rect 1111 15597 1153 15631
rect 1187 15597 1229 15631
rect 1111 15559 1229 15597
rect 1111 15525 1153 15559
rect 1187 15525 1229 15559
rect 1111 15487 1229 15525
rect 1111 15453 1153 15487
rect 1187 15453 1229 15487
rect 1111 15415 1229 15453
rect 1111 15381 1153 15415
rect 1187 15381 1229 15415
rect 1111 15332 1229 15381
rect 13761 23410 13880 23441
rect 13761 23376 13801 23410
rect 13835 23376 13880 23410
rect 13761 23338 13880 23376
rect 13761 23304 13801 23338
rect 13835 23304 13880 23338
rect 13761 23266 13880 23304
rect 13761 23232 13801 23266
rect 13835 23232 13880 23266
rect 13761 23194 13880 23232
rect 13761 23160 13801 23194
rect 13835 23160 13880 23194
rect 13761 23122 13880 23160
rect 13761 23088 13801 23122
rect 13835 23088 13880 23122
rect 13761 23050 13880 23088
rect 13761 23016 13801 23050
rect 13835 23016 13880 23050
rect 13761 22978 13880 23016
rect 13761 22944 13801 22978
rect 13835 22944 13880 22978
rect 13761 22906 13880 22944
rect 13761 22872 13801 22906
rect 13835 22872 13880 22906
rect 13761 22834 13880 22872
rect 13761 22800 13801 22834
rect 13835 22800 13880 22834
rect 13761 22762 13880 22800
rect 13761 22728 13801 22762
rect 13835 22728 13880 22762
rect 13761 22690 13880 22728
rect 13761 22656 13801 22690
rect 13835 22656 13880 22690
rect 13761 22618 13880 22656
rect 13761 22584 13801 22618
rect 13835 22584 13880 22618
rect 13761 22546 13880 22584
rect 13761 22512 13801 22546
rect 13835 22512 13880 22546
rect 13761 22474 13880 22512
rect 13761 22440 13801 22474
rect 13835 22440 13880 22474
rect 13761 22402 13880 22440
rect 13761 22368 13801 22402
rect 13835 22368 13880 22402
rect 13761 22330 13880 22368
rect 13761 22296 13801 22330
rect 13835 22296 13880 22330
rect 13761 22258 13880 22296
rect 13761 22224 13801 22258
rect 13835 22224 13880 22258
rect 13761 22186 13880 22224
rect 13761 22152 13801 22186
rect 13835 22152 13880 22186
rect 13761 22114 13880 22152
rect 13761 22080 13801 22114
rect 13835 22080 13880 22114
rect 13761 22042 13880 22080
rect 13761 22008 13801 22042
rect 13835 22008 13880 22042
rect 13761 21970 13880 22008
rect 13761 21936 13801 21970
rect 13835 21936 13880 21970
rect 13761 21898 13880 21936
rect 13761 21864 13801 21898
rect 13835 21864 13880 21898
rect 13761 21826 13880 21864
rect 13761 21792 13801 21826
rect 13835 21792 13880 21826
rect 13761 21754 13880 21792
rect 13761 21720 13801 21754
rect 13835 21720 13880 21754
rect 13761 21682 13880 21720
rect 13761 21648 13801 21682
rect 13835 21648 13880 21682
rect 13761 21610 13880 21648
rect 13761 21576 13801 21610
rect 13835 21576 13880 21610
rect 13761 21538 13880 21576
rect 13761 21504 13801 21538
rect 13835 21504 13880 21538
rect 13761 21466 13880 21504
rect 13761 21432 13801 21466
rect 13835 21432 13880 21466
rect 13761 21394 13880 21432
rect 13761 21360 13801 21394
rect 13835 21360 13880 21394
rect 13761 21322 13880 21360
rect 13761 21288 13801 21322
rect 13835 21288 13880 21322
rect 13761 21250 13880 21288
rect 13761 21216 13801 21250
rect 13835 21216 13880 21250
rect 13761 21178 13880 21216
rect 13761 21144 13801 21178
rect 13835 21144 13880 21178
rect 13761 21106 13880 21144
rect 13761 21072 13801 21106
rect 13835 21072 13880 21106
rect 13761 21034 13880 21072
rect 13761 21000 13801 21034
rect 13835 21000 13880 21034
rect 13761 20962 13880 21000
rect 13761 20928 13801 20962
rect 13835 20928 13880 20962
rect 13761 20890 13880 20928
rect 13761 20856 13801 20890
rect 13835 20856 13880 20890
rect 13761 20818 13880 20856
rect 13761 20784 13801 20818
rect 13835 20784 13880 20818
rect 13761 20746 13880 20784
rect 13761 20712 13801 20746
rect 13835 20712 13880 20746
rect 13761 20674 13880 20712
rect 13761 20640 13801 20674
rect 13835 20640 13880 20674
rect 13761 20602 13880 20640
rect 13761 20568 13801 20602
rect 13835 20568 13880 20602
rect 13761 20530 13880 20568
rect 13761 20496 13801 20530
rect 13835 20496 13880 20530
rect 13761 20458 13880 20496
rect 13761 20424 13801 20458
rect 13835 20424 13880 20458
rect 13761 20386 13880 20424
rect 13761 20352 13801 20386
rect 13835 20352 13880 20386
rect 13761 20314 13880 20352
rect 13761 20280 13801 20314
rect 13835 20280 13880 20314
rect 13761 20242 13880 20280
rect 13761 20208 13801 20242
rect 13835 20208 13880 20242
rect 13761 20170 13880 20208
rect 13761 20136 13801 20170
rect 13835 20136 13880 20170
rect 13761 20098 13880 20136
rect 13761 20064 13801 20098
rect 13835 20064 13880 20098
rect 13761 20026 13880 20064
rect 13761 19992 13801 20026
rect 13835 19992 13880 20026
rect 13761 19954 13880 19992
rect 13761 19920 13801 19954
rect 13835 19920 13880 19954
rect 13761 19882 13880 19920
rect 13761 19848 13801 19882
rect 13835 19848 13880 19882
rect 13761 19810 13880 19848
rect 13761 19776 13801 19810
rect 13835 19776 13880 19810
rect 13761 19738 13880 19776
rect 13761 19704 13801 19738
rect 13835 19704 13880 19738
rect 13761 19666 13880 19704
rect 13761 19632 13801 19666
rect 13835 19632 13880 19666
rect 13761 19594 13880 19632
rect 13761 19560 13801 19594
rect 13835 19560 13880 19594
rect 13761 19522 13880 19560
rect 13761 19488 13801 19522
rect 13835 19488 13880 19522
rect 13761 19450 13880 19488
rect 13761 19416 13801 19450
rect 13835 19416 13880 19450
rect 13761 19378 13880 19416
rect 13761 19344 13801 19378
rect 13835 19344 13880 19378
rect 13761 19306 13880 19344
rect 13761 19272 13801 19306
rect 13835 19272 13880 19306
rect 13761 19234 13880 19272
rect 13761 19200 13801 19234
rect 13835 19200 13880 19234
rect 13761 19162 13880 19200
rect 13761 19128 13801 19162
rect 13835 19128 13880 19162
rect 13761 19090 13880 19128
rect 13761 19056 13801 19090
rect 13835 19056 13880 19090
rect 13761 19018 13880 19056
rect 13761 18984 13801 19018
rect 13835 18984 13880 19018
rect 13761 18946 13880 18984
rect 13761 18912 13801 18946
rect 13835 18912 13880 18946
rect 13761 18874 13880 18912
rect 13761 18840 13801 18874
rect 13835 18840 13880 18874
rect 13761 18802 13880 18840
rect 13761 18768 13801 18802
rect 13835 18768 13880 18802
rect 13761 18730 13880 18768
rect 13761 18696 13801 18730
rect 13835 18696 13880 18730
rect 13761 18658 13880 18696
rect 13761 18624 13801 18658
rect 13835 18624 13880 18658
rect 13761 18586 13880 18624
rect 13761 18552 13801 18586
rect 13835 18552 13880 18586
rect 13761 18514 13880 18552
rect 13761 18480 13801 18514
rect 13835 18480 13880 18514
rect 13761 18442 13880 18480
rect 13761 18408 13801 18442
rect 13835 18408 13880 18442
rect 13761 18370 13880 18408
rect 13761 18336 13801 18370
rect 13835 18336 13880 18370
rect 13761 18298 13880 18336
rect 13761 18264 13801 18298
rect 13835 18264 13880 18298
rect 13761 18226 13880 18264
rect 13761 18192 13801 18226
rect 13835 18192 13880 18226
rect 13761 18154 13880 18192
rect 13761 18120 13801 18154
rect 13835 18120 13880 18154
rect 13761 18082 13880 18120
rect 13761 18048 13801 18082
rect 13835 18048 13880 18082
rect 13761 18010 13880 18048
rect 13761 17976 13801 18010
rect 13835 17976 13880 18010
rect 13761 17938 13880 17976
rect 13761 17904 13801 17938
rect 13835 17904 13880 17938
rect 13761 17866 13880 17904
rect 13761 17832 13801 17866
rect 13835 17832 13880 17866
rect 13761 17794 13880 17832
rect 13761 17760 13801 17794
rect 13835 17760 13880 17794
rect 13761 17722 13880 17760
rect 13761 17688 13801 17722
rect 13835 17688 13880 17722
rect 13761 17650 13880 17688
rect 13761 17616 13801 17650
rect 13835 17616 13880 17650
rect 13761 17578 13880 17616
rect 13761 17544 13801 17578
rect 13835 17544 13880 17578
rect 13761 17506 13880 17544
rect 13761 17472 13801 17506
rect 13835 17472 13880 17506
rect 13761 17434 13880 17472
rect 13761 17400 13801 17434
rect 13835 17400 13880 17434
rect 13761 17362 13880 17400
rect 13761 17328 13801 17362
rect 13835 17328 13880 17362
rect 13761 17290 13880 17328
rect 13761 17256 13801 17290
rect 13835 17256 13880 17290
rect 13761 17218 13880 17256
rect 13761 17184 13801 17218
rect 13835 17184 13880 17218
rect 13761 17146 13880 17184
rect 13761 17112 13801 17146
rect 13835 17112 13880 17146
rect 13761 17074 13880 17112
rect 13761 17040 13801 17074
rect 13835 17040 13880 17074
rect 13761 17002 13880 17040
rect 13761 16968 13801 17002
rect 13835 16968 13880 17002
rect 13761 16930 13880 16968
rect 13761 16896 13801 16930
rect 13835 16896 13880 16930
rect 13761 16858 13880 16896
rect 13761 16824 13801 16858
rect 13835 16824 13880 16858
rect 13761 16786 13880 16824
rect 13761 16752 13801 16786
rect 13835 16752 13880 16786
rect 13761 16714 13880 16752
rect 13761 16680 13801 16714
rect 13835 16680 13880 16714
rect 13761 16642 13880 16680
rect 13761 16608 13801 16642
rect 13835 16608 13880 16642
rect 13761 16570 13880 16608
rect 13761 16536 13801 16570
rect 13835 16536 13880 16570
rect 13761 16498 13880 16536
rect 13761 16464 13801 16498
rect 13835 16464 13880 16498
rect 13761 16426 13880 16464
rect 13761 16392 13801 16426
rect 13835 16392 13880 16426
rect 13761 16354 13880 16392
rect 13761 16320 13801 16354
rect 13835 16320 13880 16354
rect 13761 16282 13880 16320
rect 13761 16248 13801 16282
rect 13835 16248 13880 16282
rect 13761 16210 13880 16248
rect 13761 16176 13801 16210
rect 13835 16176 13880 16210
rect 13761 16138 13880 16176
rect 13761 16104 13801 16138
rect 13835 16104 13880 16138
rect 13761 16066 13880 16104
rect 13761 16032 13801 16066
rect 13835 16032 13880 16066
rect 13761 15994 13880 16032
rect 13761 15960 13801 15994
rect 13835 15960 13880 15994
rect 13761 15922 13880 15960
rect 13761 15888 13801 15922
rect 13835 15888 13880 15922
rect 13761 15850 13880 15888
rect 13761 15816 13801 15850
rect 13835 15816 13880 15850
rect 13761 15778 13880 15816
rect 13761 15744 13801 15778
rect 13835 15744 13880 15778
rect 13761 15706 13880 15744
rect 13761 15672 13801 15706
rect 13835 15672 13880 15706
rect 13761 15634 13880 15672
rect 13761 15600 13801 15634
rect 13835 15600 13880 15634
rect 13761 15562 13880 15600
rect 13761 15528 13801 15562
rect 13835 15528 13880 15562
rect 13761 15490 13880 15528
rect 13761 15456 13801 15490
rect 13835 15456 13880 15490
rect 13761 15418 13880 15456
rect 13761 15384 13801 15418
rect 13835 15384 13880 15418
rect 13761 15332 13880 15384
rect 1111 15291 13880 15332
rect 1111 15257 1290 15291
rect 1324 15257 1362 15291
rect 1396 15257 1434 15291
rect 1468 15257 1506 15291
rect 1540 15257 1578 15291
rect 1612 15257 1650 15291
rect 1684 15257 1722 15291
rect 1756 15257 1794 15291
rect 1828 15257 1866 15291
rect 1900 15257 1938 15291
rect 1972 15257 2010 15291
rect 2044 15257 2082 15291
rect 2116 15257 2154 15291
rect 2188 15257 2226 15291
rect 2260 15257 2298 15291
rect 2332 15257 2370 15291
rect 2404 15257 2442 15291
rect 2476 15257 2514 15291
rect 2548 15257 2586 15291
rect 2620 15257 2658 15291
rect 2692 15257 2730 15291
rect 2764 15257 2802 15291
rect 2836 15257 2874 15291
rect 2908 15257 2946 15291
rect 2980 15257 3018 15291
rect 3052 15257 3090 15291
rect 3124 15257 3162 15291
rect 3196 15257 3234 15291
rect 3268 15257 3306 15291
rect 3340 15257 3378 15291
rect 3412 15257 3450 15291
rect 3484 15257 3522 15291
rect 3556 15257 3594 15291
rect 3628 15257 3666 15291
rect 3700 15257 3738 15291
rect 3772 15257 3810 15291
rect 3844 15257 3882 15291
rect 3916 15257 3954 15291
rect 3988 15257 4026 15291
rect 4060 15257 4098 15291
rect 4132 15257 4170 15291
rect 4204 15257 4242 15291
rect 4276 15257 4314 15291
rect 4348 15257 4386 15291
rect 4420 15257 4458 15291
rect 4492 15257 4530 15291
rect 4564 15257 4602 15291
rect 4636 15257 4674 15291
rect 4708 15257 4746 15291
rect 4780 15257 4818 15291
rect 4852 15257 4890 15291
rect 4924 15257 4962 15291
rect 4996 15257 5034 15291
rect 5068 15257 5106 15291
rect 5140 15257 5178 15291
rect 5212 15257 5250 15291
rect 5284 15257 5322 15291
rect 5356 15257 5394 15291
rect 5428 15257 5466 15291
rect 5500 15257 5538 15291
rect 5572 15257 5610 15291
rect 5644 15257 5682 15291
rect 5716 15257 5754 15291
rect 5788 15257 5826 15291
rect 5860 15257 5898 15291
rect 5932 15257 5970 15291
rect 6004 15257 6042 15291
rect 6076 15257 6114 15291
rect 6148 15257 6186 15291
rect 6220 15257 6258 15291
rect 6292 15257 6330 15291
rect 6364 15257 6402 15291
rect 6436 15257 6474 15291
rect 6508 15257 6546 15291
rect 6580 15257 6618 15291
rect 6652 15257 6690 15291
rect 6724 15257 6762 15291
rect 6796 15257 6834 15291
rect 6868 15257 6906 15291
rect 6940 15257 6978 15291
rect 7012 15257 7050 15291
rect 7084 15257 7122 15291
rect 7156 15257 7194 15291
rect 7228 15257 7266 15291
rect 7300 15257 7338 15291
rect 7372 15257 7410 15291
rect 7444 15257 7482 15291
rect 7516 15257 7554 15291
rect 7588 15257 7626 15291
rect 7660 15257 7698 15291
rect 7732 15257 7770 15291
rect 7804 15257 7842 15291
rect 7876 15257 7914 15291
rect 7948 15257 7986 15291
rect 8020 15257 8058 15291
rect 8092 15257 8130 15291
rect 8164 15257 8202 15291
rect 8236 15257 8274 15291
rect 8308 15257 8346 15291
rect 8380 15257 8418 15291
rect 8452 15257 8490 15291
rect 8524 15257 8562 15291
rect 8596 15257 8634 15291
rect 8668 15257 8706 15291
rect 8740 15257 8778 15291
rect 8812 15257 8850 15291
rect 8884 15257 8922 15291
rect 8956 15257 8994 15291
rect 9028 15257 9066 15291
rect 9100 15257 9138 15291
rect 9172 15257 9210 15291
rect 9244 15257 9282 15291
rect 9316 15257 9354 15291
rect 9388 15257 9426 15291
rect 9460 15257 9498 15291
rect 9532 15257 9570 15291
rect 9604 15257 9642 15291
rect 9676 15257 9714 15291
rect 9748 15257 9786 15291
rect 9820 15257 9858 15291
rect 9892 15257 9930 15291
rect 9964 15257 10002 15291
rect 10036 15257 10074 15291
rect 10108 15257 10146 15291
rect 10180 15257 10218 15291
rect 10252 15257 10290 15291
rect 10324 15257 10362 15291
rect 10396 15257 10434 15291
rect 10468 15257 10506 15291
rect 10540 15257 10578 15291
rect 10612 15257 10650 15291
rect 10684 15257 10722 15291
rect 10756 15257 10794 15291
rect 10828 15257 10866 15291
rect 10900 15257 10938 15291
rect 10972 15257 11010 15291
rect 11044 15257 11082 15291
rect 11116 15257 11154 15291
rect 11188 15257 11226 15291
rect 11260 15257 11298 15291
rect 11332 15257 11370 15291
rect 11404 15257 11442 15291
rect 11476 15257 11514 15291
rect 11548 15257 11586 15291
rect 11620 15257 11658 15291
rect 11692 15257 11730 15291
rect 11764 15257 11802 15291
rect 11836 15257 11874 15291
rect 11908 15257 11946 15291
rect 11980 15257 12018 15291
rect 12052 15257 12090 15291
rect 12124 15257 12162 15291
rect 12196 15257 12234 15291
rect 12268 15257 12306 15291
rect 12340 15257 12378 15291
rect 12412 15257 12450 15291
rect 12484 15257 12522 15291
rect 12556 15257 12594 15291
rect 12628 15257 12666 15291
rect 12700 15257 12738 15291
rect 12772 15257 12810 15291
rect 12844 15257 12882 15291
rect 12916 15257 12954 15291
rect 12988 15257 13026 15291
rect 13060 15257 13098 15291
rect 13132 15257 13170 15291
rect 13204 15257 13242 15291
rect 13276 15257 13314 15291
rect 13348 15257 13386 15291
rect 13420 15257 13458 15291
rect 13492 15257 13530 15291
rect 13564 15257 13602 15291
rect 13636 15257 13674 15291
rect 13708 15257 13880 15291
rect 1111 15214 13880 15257
rect 14091 23416 14114 23450
rect 14148 23416 14211 23450
rect 14091 23378 14211 23416
rect 14091 23344 14114 23378
rect 14148 23344 14211 23378
rect 14091 23306 14211 23344
rect 14091 23272 14114 23306
rect 14148 23272 14211 23306
rect 14091 23234 14211 23272
rect 14091 23200 14114 23234
rect 14148 23200 14211 23234
rect 14091 23162 14211 23200
rect 14091 23128 14114 23162
rect 14148 23128 14211 23162
rect 14091 23090 14211 23128
rect 14091 23056 14114 23090
rect 14148 23056 14211 23090
rect 14091 23018 14211 23056
rect 14091 22984 14114 23018
rect 14148 22984 14211 23018
rect 14091 22946 14211 22984
rect 14091 22912 14114 22946
rect 14148 22912 14211 22946
rect 14091 22874 14211 22912
rect 14091 22840 14114 22874
rect 14148 22840 14211 22874
rect 14091 22802 14211 22840
rect 14091 22768 14114 22802
rect 14148 22768 14211 22802
rect 14091 22730 14211 22768
rect 14091 22696 14114 22730
rect 14148 22696 14211 22730
rect 14091 22658 14211 22696
rect 14091 22624 14114 22658
rect 14148 22624 14211 22658
rect 14091 22586 14211 22624
rect 14091 22552 14114 22586
rect 14148 22552 14211 22586
rect 14091 22514 14211 22552
rect 14091 22480 14114 22514
rect 14148 22480 14211 22514
rect 14091 22442 14211 22480
rect 14091 22408 14114 22442
rect 14148 22408 14211 22442
rect 14091 22370 14211 22408
rect 14091 22336 14114 22370
rect 14148 22336 14211 22370
rect 14091 22298 14211 22336
rect 14091 22264 14114 22298
rect 14148 22264 14211 22298
rect 14091 22226 14211 22264
rect 14091 22192 14114 22226
rect 14148 22192 14211 22226
rect 14091 22154 14211 22192
rect 14091 22120 14114 22154
rect 14148 22120 14211 22154
rect 14091 22082 14211 22120
rect 14091 22048 14114 22082
rect 14148 22048 14211 22082
rect 14091 22010 14211 22048
rect 14091 21976 14114 22010
rect 14148 21976 14211 22010
rect 14091 21938 14211 21976
rect 14091 21904 14114 21938
rect 14148 21904 14211 21938
rect 14091 21866 14211 21904
rect 14091 21832 14114 21866
rect 14148 21832 14211 21866
rect 14091 21794 14211 21832
rect 14091 21760 14114 21794
rect 14148 21760 14211 21794
rect 14091 21722 14211 21760
rect 14091 21688 14114 21722
rect 14148 21688 14211 21722
rect 14091 21650 14211 21688
rect 14091 21616 14114 21650
rect 14148 21616 14211 21650
rect 14091 21578 14211 21616
rect 14091 21544 14114 21578
rect 14148 21544 14211 21578
rect 14091 21506 14211 21544
rect 14091 21472 14114 21506
rect 14148 21472 14211 21506
rect 14091 21434 14211 21472
rect 14091 21400 14114 21434
rect 14148 21400 14211 21434
rect 14091 21362 14211 21400
rect 14091 21328 14114 21362
rect 14148 21328 14211 21362
rect 14091 21290 14211 21328
rect 14091 21256 14114 21290
rect 14148 21256 14211 21290
rect 14091 21218 14211 21256
rect 14091 21184 14114 21218
rect 14148 21184 14211 21218
rect 14091 21146 14211 21184
rect 14091 21112 14114 21146
rect 14148 21112 14211 21146
rect 14091 21074 14211 21112
rect 14091 21040 14114 21074
rect 14148 21040 14211 21074
rect 14091 21002 14211 21040
rect 14091 20968 14114 21002
rect 14148 20968 14211 21002
rect 14091 20930 14211 20968
rect 14091 20896 14114 20930
rect 14148 20896 14211 20930
rect 14091 20858 14211 20896
rect 14091 20824 14114 20858
rect 14148 20824 14211 20858
rect 14091 20786 14211 20824
rect 14091 20752 14114 20786
rect 14148 20752 14211 20786
rect 14091 20714 14211 20752
rect 14091 20680 14114 20714
rect 14148 20680 14211 20714
rect 14091 20642 14211 20680
rect 14091 20608 14114 20642
rect 14148 20608 14211 20642
rect 14091 20570 14211 20608
rect 14091 20536 14114 20570
rect 14148 20536 14211 20570
rect 14091 20498 14211 20536
rect 14091 20464 14114 20498
rect 14148 20464 14211 20498
rect 14091 20426 14211 20464
rect 14091 20392 14114 20426
rect 14148 20392 14211 20426
rect 14091 20354 14211 20392
rect 14091 20320 14114 20354
rect 14148 20320 14211 20354
rect 14091 20282 14211 20320
rect 14091 20248 14114 20282
rect 14148 20248 14211 20282
rect 14091 20210 14211 20248
rect 14091 20176 14114 20210
rect 14148 20176 14211 20210
rect 14091 20138 14211 20176
rect 14091 20104 14114 20138
rect 14148 20104 14211 20138
rect 14091 20066 14211 20104
rect 14091 20032 14114 20066
rect 14148 20032 14211 20066
rect 14091 19994 14211 20032
rect 14091 19960 14114 19994
rect 14148 19960 14211 19994
rect 14091 19922 14211 19960
rect 14091 19888 14114 19922
rect 14148 19888 14211 19922
rect 14091 19850 14211 19888
rect 14091 19816 14114 19850
rect 14148 19816 14211 19850
rect 14091 19778 14211 19816
rect 14091 19744 14114 19778
rect 14148 19744 14211 19778
rect 14091 19706 14211 19744
rect 14091 19672 14114 19706
rect 14148 19672 14211 19706
rect 14091 19634 14211 19672
rect 14091 19600 14114 19634
rect 14148 19600 14211 19634
rect 14091 19562 14211 19600
rect 14091 19528 14114 19562
rect 14148 19528 14211 19562
rect 14091 19490 14211 19528
rect 14091 19456 14114 19490
rect 14148 19456 14211 19490
rect 14091 19418 14211 19456
rect 14091 19384 14114 19418
rect 14148 19384 14211 19418
rect 14091 19346 14211 19384
rect 14091 19312 14114 19346
rect 14148 19312 14211 19346
rect 14091 19274 14211 19312
rect 14091 19240 14114 19274
rect 14148 19240 14211 19274
rect 14091 19202 14211 19240
rect 14091 19168 14114 19202
rect 14148 19168 14211 19202
rect 14091 19130 14211 19168
rect 14091 19096 14114 19130
rect 14148 19096 14211 19130
rect 14091 19058 14211 19096
rect 14091 19024 14114 19058
rect 14148 19024 14211 19058
rect 14091 18986 14211 19024
rect 14091 18952 14114 18986
rect 14148 18952 14211 18986
rect 14091 18914 14211 18952
rect 14091 18880 14114 18914
rect 14148 18880 14211 18914
rect 14091 18842 14211 18880
rect 14091 18808 14114 18842
rect 14148 18808 14211 18842
rect 14091 18770 14211 18808
rect 14091 18736 14114 18770
rect 14148 18736 14211 18770
rect 14091 18698 14211 18736
rect 14091 18664 14114 18698
rect 14148 18664 14211 18698
rect 14091 18626 14211 18664
rect 14091 18592 14114 18626
rect 14148 18592 14211 18626
rect 14091 18554 14211 18592
rect 14091 18520 14114 18554
rect 14148 18520 14211 18554
rect 14091 18482 14211 18520
rect 14091 18448 14114 18482
rect 14148 18448 14211 18482
rect 14091 18410 14211 18448
rect 14091 18376 14114 18410
rect 14148 18376 14211 18410
rect 14091 18338 14211 18376
rect 14091 18304 14114 18338
rect 14148 18304 14211 18338
rect 14091 18266 14211 18304
rect 14091 18232 14114 18266
rect 14148 18232 14211 18266
rect 14091 18194 14211 18232
rect 14091 18160 14114 18194
rect 14148 18160 14211 18194
rect 14091 18122 14211 18160
rect 14091 18088 14114 18122
rect 14148 18088 14211 18122
rect 14091 18050 14211 18088
rect 14091 18016 14114 18050
rect 14148 18016 14211 18050
rect 14091 17978 14211 18016
rect 14091 17944 14114 17978
rect 14148 17944 14211 17978
rect 14091 17906 14211 17944
rect 14091 17872 14114 17906
rect 14148 17872 14211 17906
rect 14091 17834 14211 17872
rect 14091 17800 14114 17834
rect 14148 17800 14211 17834
rect 14091 17762 14211 17800
rect 14091 17728 14114 17762
rect 14148 17728 14211 17762
rect 14091 17690 14211 17728
rect 14091 17656 14114 17690
rect 14148 17656 14211 17690
rect 14091 17618 14211 17656
rect 14091 17584 14114 17618
rect 14148 17584 14211 17618
rect 14091 17546 14211 17584
rect 14091 17512 14114 17546
rect 14148 17512 14211 17546
rect 14091 17474 14211 17512
rect 14091 17440 14114 17474
rect 14148 17440 14211 17474
rect 14091 17402 14211 17440
rect 14091 17368 14114 17402
rect 14148 17368 14211 17402
rect 14091 17330 14211 17368
rect 14091 17296 14114 17330
rect 14148 17296 14211 17330
rect 14091 17258 14211 17296
rect 14091 17224 14114 17258
rect 14148 17224 14211 17258
rect 14091 17186 14211 17224
rect 14091 17152 14114 17186
rect 14148 17152 14211 17186
rect 14091 17114 14211 17152
rect 14091 17080 14114 17114
rect 14148 17080 14211 17114
rect 14091 17042 14211 17080
rect 14091 17008 14114 17042
rect 14148 17008 14211 17042
rect 14091 16970 14211 17008
rect 14091 16936 14114 16970
rect 14148 16936 14211 16970
rect 14091 16898 14211 16936
rect 14091 16864 14114 16898
rect 14148 16864 14211 16898
rect 14091 16826 14211 16864
rect 14091 16792 14114 16826
rect 14148 16792 14211 16826
rect 14091 16754 14211 16792
rect 14091 16720 14114 16754
rect 14148 16720 14211 16754
rect 14091 16682 14211 16720
rect 14091 16648 14114 16682
rect 14148 16648 14211 16682
rect 14091 16610 14211 16648
rect 14091 16576 14114 16610
rect 14148 16576 14211 16610
rect 14091 16538 14211 16576
rect 14091 16504 14114 16538
rect 14148 16504 14211 16538
rect 14091 16466 14211 16504
rect 14091 16432 14114 16466
rect 14148 16432 14211 16466
rect 14091 16394 14211 16432
rect 14091 16360 14114 16394
rect 14148 16360 14211 16394
rect 14091 16322 14211 16360
rect 14091 16288 14114 16322
rect 14148 16288 14211 16322
rect 14091 16250 14211 16288
rect 14091 16216 14114 16250
rect 14148 16216 14211 16250
rect 14091 16178 14211 16216
rect 14091 16144 14114 16178
rect 14148 16144 14211 16178
rect 14091 16106 14211 16144
rect 14091 16072 14114 16106
rect 14148 16072 14211 16106
rect 14091 16034 14211 16072
rect 14091 16000 14114 16034
rect 14148 16000 14211 16034
rect 14091 15962 14211 16000
rect 14091 15928 14114 15962
rect 14148 15928 14211 15962
rect 14091 15890 14211 15928
rect 14091 15856 14114 15890
rect 14148 15856 14211 15890
rect 14091 15818 14211 15856
rect 14091 15784 14114 15818
rect 14148 15784 14211 15818
rect 14091 15746 14211 15784
rect 14091 15712 14114 15746
rect 14148 15712 14211 15746
rect 14091 15674 14211 15712
rect 14091 15640 14114 15674
rect 14148 15640 14211 15674
rect 14091 15602 14211 15640
rect 14091 15568 14114 15602
rect 14148 15568 14211 15602
rect 14091 15530 14211 15568
rect 14091 15496 14114 15530
rect 14148 15496 14211 15530
rect 14091 15458 14211 15496
rect 14091 15424 14114 15458
rect 14148 15424 14211 15458
rect 14091 15386 14211 15424
rect 14091 15352 14114 15386
rect 14148 15352 14211 15386
rect 14091 15314 14211 15352
rect 14091 15280 14114 15314
rect 14148 15280 14211 15314
rect 14091 15242 14211 15280
rect 749 15143 799 15177
rect 833 15143 869 15177
rect 749 15105 869 15143
rect 749 15071 799 15105
rect 833 15071 869 15105
rect 749 14976 869 15071
rect 14091 15208 14114 15242
rect 14148 15208 14211 15242
rect 14091 15170 14211 15208
rect 14091 15136 14114 15170
rect 14148 15136 14211 15170
rect 14091 15098 14211 15136
rect 14091 15064 14114 15098
rect 14148 15064 14211 15098
tri 869 14976 909 15016 sw
tri 14051 14976 14091 15016 se
rect 14091 14976 14211 15064
rect 749 14956 14211 14976
tri 749 14856 849 14956 ne
rect 849 14955 14111 14956
rect 849 14921 883 14955
rect 917 14921 955 14955
rect 989 14921 1027 14955
rect 1061 14921 1099 14955
rect 1133 14921 1171 14955
rect 1205 14921 1243 14955
rect 1277 14921 1315 14955
rect 1349 14921 1387 14955
rect 1421 14921 1459 14955
rect 1493 14921 1531 14955
rect 1565 14921 1603 14955
rect 1637 14921 1675 14955
rect 1709 14921 1747 14955
rect 1781 14921 1819 14955
rect 1853 14921 1891 14955
rect 1925 14921 1963 14955
rect 1997 14921 2035 14955
rect 2069 14921 2107 14955
rect 2141 14921 2179 14955
rect 2213 14921 2251 14955
rect 2285 14921 2323 14955
rect 2357 14921 2395 14955
rect 2429 14921 2467 14955
rect 2501 14921 2539 14955
rect 2573 14921 2611 14955
rect 2645 14921 2683 14955
rect 2717 14921 2755 14955
rect 2789 14921 2827 14955
rect 2861 14921 2899 14955
rect 2933 14921 2971 14955
rect 3005 14921 3043 14955
rect 3077 14921 3115 14955
rect 3149 14921 3187 14955
rect 3221 14921 3259 14955
rect 3293 14921 3331 14955
rect 3365 14921 3403 14955
rect 3437 14921 3475 14955
rect 3509 14921 3547 14955
rect 3581 14921 3619 14955
rect 3653 14921 3691 14955
rect 3725 14921 3763 14955
rect 3797 14921 3835 14955
rect 3869 14921 3907 14955
rect 3941 14921 3979 14955
rect 4013 14921 4051 14955
rect 4085 14921 4123 14955
rect 4157 14921 4195 14955
rect 4229 14921 4267 14955
rect 4301 14921 4339 14955
rect 4373 14921 4411 14955
rect 4445 14921 4483 14955
rect 4517 14921 4555 14955
rect 4589 14921 4627 14955
rect 4661 14921 4699 14955
rect 4733 14921 4771 14955
rect 4805 14921 4843 14955
rect 4877 14921 4915 14955
rect 4949 14921 4987 14955
rect 5021 14921 5059 14955
rect 5093 14921 5131 14955
rect 5165 14921 5203 14955
rect 5237 14921 5275 14955
rect 5309 14921 5347 14955
rect 5381 14921 5419 14955
rect 5453 14921 5491 14955
rect 5525 14921 5563 14955
rect 5597 14921 5635 14955
rect 5669 14921 5707 14955
rect 5741 14921 5779 14955
rect 5813 14921 5851 14955
rect 5885 14921 5923 14955
rect 5957 14921 5995 14955
rect 6029 14921 6067 14955
rect 6101 14921 6139 14955
rect 6173 14921 6211 14955
rect 6245 14921 6283 14955
rect 6317 14921 6355 14955
rect 6389 14921 6427 14955
rect 6461 14921 6499 14955
rect 6533 14921 6571 14955
rect 6605 14921 6643 14955
rect 6677 14921 6715 14955
rect 6749 14921 6787 14955
rect 6821 14921 6859 14955
rect 6893 14921 6931 14955
rect 6965 14921 7003 14955
rect 7037 14921 7075 14955
rect 7109 14921 7147 14955
rect 7181 14921 7219 14955
rect 7253 14921 7291 14955
rect 7325 14921 7363 14955
rect 7397 14921 7435 14955
rect 7469 14921 7507 14955
rect 7541 14921 7579 14955
rect 7613 14921 7651 14955
rect 7685 14921 7723 14955
rect 7757 14921 7795 14955
rect 7829 14921 7867 14955
rect 7901 14921 7939 14955
rect 7973 14921 8011 14955
rect 8045 14921 8083 14955
rect 8117 14921 8155 14955
rect 8189 14921 8227 14955
rect 8261 14921 8299 14955
rect 8333 14921 8371 14955
rect 8405 14921 8443 14955
rect 8477 14921 8515 14955
rect 8549 14921 8587 14955
rect 8621 14921 8659 14955
rect 8693 14921 8731 14955
rect 8765 14921 8803 14955
rect 8837 14921 8875 14955
rect 8909 14921 8947 14955
rect 8981 14921 9019 14955
rect 9053 14921 9091 14955
rect 9125 14921 9163 14955
rect 9197 14921 9235 14955
rect 9269 14921 9307 14955
rect 9341 14921 9379 14955
rect 9413 14921 9451 14955
rect 9485 14921 9523 14955
rect 9557 14921 9595 14955
rect 9629 14921 9667 14955
rect 9701 14921 9739 14955
rect 9773 14921 9811 14955
rect 9845 14921 9883 14955
rect 9917 14921 9955 14955
rect 9989 14921 10027 14955
rect 10061 14921 10099 14955
rect 10133 14921 10171 14955
rect 10205 14921 10243 14955
rect 10277 14921 10315 14955
rect 10349 14921 10387 14955
rect 10421 14921 10459 14955
rect 10493 14921 10531 14955
rect 10565 14921 10603 14955
rect 10637 14921 10675 14955
rect 10709 14921 10747 14955
rect 10781 14921 10819 14955
rect 10853 14921 10891 14955
rect 10925 14921 10963 14955
rect 10997 14921 11035 14955
rect 11069 14921 11107 14955
rect 11141 14921 11179 14955
rect 11213 14921 11251 14955
rect 11285 14921 11323 14955
rect 11357 14921 11395 14955
rect 11429 14921 11467 14955
rect 11501 14921 11539 14955
rect 11573 14921 11611 14955
rect 11645 14921 11683 14955
rect 11717 14921 11755 14955
rect 11789 14921 11827 14955
rect 11861 14921 11899 14955
rect 11933 14921 11971 14955
rect 12005 14921 12043 14955
rect 12077 14921 12115 14955
rect 12149 14921 12187 14955
rect 12221 14921 12259 14955
rect 12293 14921 12331 14955
rect 12365 14921 12403 14955
rect 12437 14921 12475 14955
rect 12509 14921 12547 14955
rect 12581 14921 12619 14955
rect 12653 14921 12691 14955
rect 12725 14921 12763 14955
rect 12797 14921 12835 14955
rect 12869 14921 12907 14955
rect 12941 14921 12979 14955
rect 13013 14921 13051 14955
rect 13085 14921 13123 14955
rect 13157 14921 13195 14955
rect 13229 14921 13267 14955
rect 13301 14921 13339 14955
rect 13373 14921 13411 14955
rect 13445 14921 13483 14955
rect 13517 14921 13555 14955
rect 13589 14921 13627 14955
rect 13661 14921 13699 14955
rect 13733 14921 13771 14955
rect 13805 14921 13843 14955
rect 13877 14921 13915 14955
rect 13949 14921 13987 14955
rect 14021 14921 14111 14955
rect 849 14856 14111 14921
tri 14111 14856 14211 14956 nw
rect 14531 36041 14606 36075
rect 14640 36041 14716 36075
rect 14531 36003 14716 36041
rect 14531 35969 14606 36003
rect 14640 35969 14716 36003
rect 14531 35931 14716 35969
rect 14531 35897 14606 35931
rect 14640 35897 14716 35931
rect 14531 35859 14716 35897
rect 14531 35825 14606 35859
rect 14640 35825 14716 35859
rect 14531 35787 14716 35825
rect 14531 35753 14606 35787
rect 14640 35753 14716 35787
rect 14531 35715 14716 35753
rect 14531 35681 14606 35715
rect 14640 35681 14716 35715
rect 14531 35643 14716 35681
rect 14531 35609 14606 35643
rect 14640 35609 14716 35643
rect 14531 35571 14716 35609
rect 14531 35537 14606 35571
rect 14640 35537 14716 35571
rect 14531 35499 14716 35537
rect 14531 35465 14606 35499
rect 14640 35465 14716 35499
rect 14531 35427 14716 35465
rect 14531 35393 14606 35427
rect 14640 35393 14716 35427
rect 14531 35355 14716 35393
rect 14531 35321 14606 35355
rect 14640 35321 14716 35355
rect 14531 35283 14716 35321
rect 14531 35249 14606 35283
rect 14640 35249 14716 35283
rect 14531 35211 14716 35249
rect 14531 35177 14606 35211
rect 14640 35177 14716 35211
rect 14531 35139 14716 35177
rect 14531 35105 14606 35139
rect 14640 35105 14716 35139
rect 14531 35067 14716 35105
rect 14531 35033 14606 35067
rect 14640 35033 14716 35067
rect 14531 34995 14716 35033
rect 14531 34961 14606 34995
rect 14640 34961 14716 34995
rect 14531 34923 14716 34961
rect 14531 34889 14606 34923
rect 14640 34889 14716 34923
rect 14531 34851 14716 34889
rect 14531 34817 14606 34851
rect 14640 34817 14716 34851
rect 14531 34779 14716 34817
rect 14531 34745 14606 34779
rect 14640 34745 14716 34779
rect 14531 34707 14716 34745
rect 14531 34673 14606 34707
rect 14640 34673 14716 34707
rect 14531 34635 14716 34673
rect 14531 34601 14606 34635
rect 14640 34601 14716 34635
rect 14531 34563 14716 34601
rect 14531 34529 14606 34563
rect 14640 34529 14716 34563
rect 14531 34491 14716 34529
rect 14531 34457 14606 34491
rect 14640 34457 14716 34491
rect 14531 34419 14716 34457
rect 14531 34385 14606 34419
rect 14640 34385 14716 34419
rect 14531 34347 14716 34385
rect 14531 34313 14606 34347
rect 14640 34313 14716 34347
rect 14531 34275 14716 34313
rect 14531 34241 14606 34275
rect 14640 34241 14716 34275
rect 14531 34203 14716 34241
rect 14531 34169 14606 34203
rect 14640 34169 14716 34203
rect 14531 34131 14716 34169
rect 14531 34097 14606 34131
rect 14640 34097 14716 34131
rect 14531 34059 14716 34097
rect 14531 34025 14606 34059
rect 14640 34025 14716 34059
rect 14531 33987 14716 34025
rect 14531 33953 14606 33987
rect 14640 33953 14716 33987
rect 14531 33915 14716 33953
rect 14531 33881 14606 33915
rect 14640 33881 14716 33915
rect 14531 33843 14716 33881
rect 14531 33809 14606 33843
rect 14640 33809 14716 33843
rect 14531 33771 14716 33809
rect 14531 33737 14606 33771
rect 14640 33737 14716 33771
rect 14531 33699 14716 33737
rect 14531 33665 14606 33699
rect 14640 33665 14716 33699
rect 14531 33627 14716 33665
rect 14531 33593 14606 33627
rect 14640 33593 14716 33627
rect 14531 33555 14716 33593
rect 14531 33521 14606 33555
rect 14640 33521 14716 33555
rect 14531 33483 14716 33521
rect 14531 33449 14606 33483
rect 14640 33449 14716 33483
rect 14531 33411 14716 33449
rect 14531 33377 14606 33411
rect 14640 33377 14716 33411
rect 14531 33339 14716 33377
rect 14531 33305 14606 33339
rect 14640 33305 14716 33339
rect 14531 33267 14716 33305
rect 14531 33233 14606 33267
rect 14640 33233 14716 33267
rect 14531 33195 14716 33233
rect 14531 33161 14606 33195
rect 14640 33161 14716 33195
rect 14531 33123 14716 33161
rect 14531 33089 14606 33123
rect 14640 33089 14716 33123
rect 14531 33051 14716 33089
rect 14531 33017 14606 33051
rect 14640 33017 14716 33051
rect 14531 32979 14716 33017
rect 14531 32945 14606 32979
rect 14640 32945 14716 32979
rect 14531 32907 14716 32945
rect 14531 32873 14606 32907
rect 14640 32873 14716 32907
rect 14531 32835 14716 32873
rect 14531 32801 14606 32835
rect 14640 32801 14716 32835
rect 14531 32763 14716 32801
rect 14531 32729 14606 32763
rect 14640 32729 14716 32763
rect 14531 32691 14716 32729
rect 14531 32657 14606 32691
rect 14640 32657 14716 32691
rect 14531 32619 14716 32657
rect 14531 32585 14606 32619
rect 14640 32585 14716 32619
rect 14531 32547 14716 32585
rect 14531 32513 14606 32547
rect 14640 32513 14716 32547
rect 14531 32475 14716 32513
rect 14531 32441 14606 32475
rect 14640 32441 14716 32475
rect 14531 32403 14716 32441
rect 14531 32369 14606 32403
rect 14640 32369 14716 32403
rect 14531 32331 14716 32369
rect 14531 32297 14606 32331
rect 14640 32297 14716 32331
rect 14531 32259 14716 32297
rect 14531 32225 14606 32259
rect 14640 32225 14716 32259
rect 14531 32187 14716 32225
rect 14531 32153 14606 32187
rect 14640 32153 14716 32187
rect 14531 32115 14716 32153
rect 14531 32081 14606 32115
rect 14640 32081 14716 32115
rect 14531 32043 14716 32081
rect 14531 32009 14606 32043
rect 14640 32009 14716 32043
rect 14531 31971 14716 32009
rect 14531 31937 14606 31971
rect 14640 31937 14716 31971
rect 14531 31899 14716 31937
rect 14531 31865 14606 31899
rect 14640 31865 14716 31899
rect 14531 31827 14716 31865
rect 14531 31793 14606 31827
rect 14640 31793 14716 31827
rect 14531 31755 14716 31793
rect 14531 31721 14606 31755
rect 14640 31721 14716 31755
rect 14531 31683 14716 31721
rect 14531 31649 14606 31683
rect 14640 31649 14716 31683
rect 14531 31611 14716 31649
rect 14531 31577 14606 31611
rect 14640 31577 14716 31611
rect 14531 31539 14716 31577
rect 14531 31505 14606 31539
rect 14640 31505 14716 31539
rect 14531 31467 14716 31505
rect 14531 31433 14606 31467
rect 14640 31433 14716 31467
rect 14531 31395 14716 31433
rect 14531 31361 14606 31395
rect 14640 31361 14716 31395
rect 14531 31323 14716 31361
rect 14531 31289 14606 31323
rect 14640 31289 14716 31323
rect 14531 31251 14716 31289
rect 14531 31217 14606 31251
rect 14640 31217 14716 31251
rect 14531 31179 14716 31217
rect 14531 31145 14606 31179
rect 14640 31145 14716 31179
rect 14531 31107 14716 31145
rect 14531 31073 14606 31107
rect 14640 31073 14716 31107
rect 14531 31035 14716 31073
rect 14531 31001 14606 31035
rect 14640 31001 14716 31035
rect 14531 30963 14716 31001
rect 14531 30929 14606 30963
rect 14640 30929 14716 30963
rect 14531 30891 14716 30929
rect 14531 30857 14606 30891
rect 14640 30857 14716 30891
rect 14531 30819 14716 30857
rect 14531 30785 14606 30819
rect 14640 30785 14716 30819
rect 14531 30747 14716 30785
rect 14531 30713 14606 30747
rect 14640 30713 14716 30747
rect 14531 30675 14716 30713
rect 14531 30641 14606 30675
rect 14640 30641 14716 30675
rect 14531 30603 14716 30641
rect 14531 30569 14606 30603
rect 14640 30569 14716 30603
rect 14531 30531 14716 30569
rect 14531 30497 14606 30531
rect 14640 30497 14716 30531
rect 14531 30459 14716 30497
rect 14531 30425 14606 30459
rect 14640 30425 14716 30459
rect 14531 30387 14716 30425
rect 14531 30353 14606 30387
rect 14640 30353 14716 30387
rect 14531 30315 14716 30353
rect 14531 30281 14606 30315
rect 14640 30281 14716 30315
rect 14531 30243 14716 30281
rect 14531 30209 14606 30243
rect 14640 30209 14716 30243
rect 14531 30171 14716 30209
rect 14531 30137 14606 30171
rect 14640 30137 14716 30171
rect 14531 30099 14716 30137
rect 14531 30065 14606 30099
rect 14640 30065 14716 30099
rect 14531 30027 14716 30065
rect 14531 29993 14606 30027
rect 14640 29993 14716 30027
rect 14531 29955 14716 29993
rect 14531 29921 14606 29955
rect 14640 29921 14716 29955
rect 14531 29883 14716 29921
rect 14531 29849 14606 29883
rect 14640 29849 14716 29883
rect 14531 29811 14716 29849
rect 14531 29777 14606 29811
rect 14640 29777 14716 29811
rect 14531 29739 14716 29777
rect 14531 29705 14606 29739
rect 14640 29705 14716 29739
rect 14531 29667 14716 29705
rect 14531 29633 14606 29667
rect 14640 29633 14716 29667
rect 14531 29595 14716 29633
rect 14531 29561 14606 29595
rect 14640 29561 14716 29595
rect 14531 29523 14716 29561
rect 14531 29489 14606 29523
rect 14640 29489 14716 29523
rect 14531 29451 14716 29489
rect 14531 29417 14606 29451
rect 14640 29417 14716 29451
rect 14531 29379 14716 29417
rect 14531 29345 14606 29379
rect 14640 29345 14716 29379
rect 14531 29307 14716 29345
rect 14531 29273 14606 29307
rect 14640 29273 14716 29307
rect 14531 29235 14716 29273
rect 14531 29201 14606 29235
rect 14640 29201 14716 29235
rect 14531 29163 14716 29201
rect 14531 29129 14606 29163
rect 14640 29129 14716 29163
rect 14531 29091 14716 29129
rect 14531 29057 14606 29091
rect 14640 29057 14716 29091
rect 14531 29019 14716 29057
rect 14531 28985 14606 29019
rect 14640 28985 14716 29019
rect 14531 28947 14716 28985
rect 14531 28913 14606 28947
rect 14640 28913 14716 28947
rect 14531 28875 14716 28913
rect 14531 28841 14606 28875
rect 14640 28841 14716 28875
rect 14531 28803 14716 28841
rect 14531 28769 14606 28803
rect 14640 28769 14716 28803
rect 14531 28731 14716 28769
rect 14531 28697 14606 28731
rect 14640 28697 14716 28731
rect 14531 28659 14716 28697
rect 14531 28625 14606 28659
rect 14640 28625 14716 28659
rect 14531 28587 14716 28625
rect 14531 28553 14606 28587
rect 14640 28553 14716 28587
rect 14531 28515 14716 28553
rect 14531 28481 14606 28515
rect 14640 28481 14716 28515
rect 14531 28443 14716 28481
rect 14531 28409 14606 28443
rect 14640 28409 14716 28443
rect 14531 28371 14716 28409
rect 14531 28337 14606 28371
rect 14640 28337 14716 28371
rect 14531 28299 14716 28337
rect 14531 28265 14606 28299
rect 14640 28265 14716 28299
rect 14531 28227 14716 28265
rect 14531 28193 14606 28227
rect 14640 28193 14716 28227
rect 14531 28155 14716 28193
rect 14531 28121 14606 28155
rect 14640 28121 14716 28155
rect 14531 28083 14716 28121
rect 14531 28049 14606 28083
rect 14640 28049 14716 28083
rect 14531 28011 14716 28049
rect 14531 27977 14606 28011
rect 14640 27977 14716 28011
rect 14531 27939 14716 27977
rect 14531 27905 14606 27939
rect 14640 27905 14716 27939
rect 14531 27867 14716 27905
rect 14531 27833 14606 27867
rect 14640 27833 14716 27867
rect 14531 27795 14716 27833
rect 14531 27761 14606 27795
rect 14640 27761 14716 27795
rect 14531 27723 14716 27761
rect 14531 27689 14606 27723
rect 14640 27689 14716 27723
rect 14531 27651 14716 27689
rect 14531 27617 14606 27651
rect 14640 27617 14716 27651
rect 14531 27579 14716 27617
rect 14531 27545 14606 27579
rect 14640 27545 14716 27579
rect 14531 27507 14716 27545
rect 14531 27473 14606 27507
rect 14640 27473 14716 27507
rect 14531 27435 14716 27473
rect 14531 27401 14606 27435
rect 14640 27401 14716 27435
rect 14531 27363 14716 27401
rect 14531 27329 14606 27363
rect 14640 27329 14716 27363
rect 14531 27291 14716 27329
rect 14531 27257 14606 27291
rect 14640 27257 14716 27291
rect 14531 27219 14716 27257
rect 14531 27185 14606 27219
rect 14640 27185 14716 27219
rect 14531 27147 14716 27185
rect 14531 27113 14606 27147
rect 14640 27113 14716 27147
rect 14531 27075 14716 27113
rect 14531 27041 14606 27075
rect 14640 27041 14716 27075
rect 14531 27003 14716 27041
rect 14531 26969 14606 27003
rect 14640 26969 14716 27003
rect 14531 26931 14716 26969
rect 14531 26897 14606 26931
rect 14640 26897 14716 26931
rect 14531 26859 14716 26897
rect 14531 26825 14606 26859
rect 14640 26825 14716 26859
rect 14531 26787 14716 26825
rect 14531 26753 14606 26787
rect 14640 26753 14716 26787
rect 14531 26715 14716 26753
rect 14531 26681 14606 26715
rect 14640 26681 14716 26715
rect 14531 26643 14716 26681
rect 14531 26609 14606 26643
rect 14640 26609 14716 26643
rect 14531 26571 14716 26609
rect 14531 26537 14606 26571
rect 14640 26537 14716 26571
rect 14531 26499 14716 26537
rect 14531 26465 14606 26499
rect 14640 26465 14716 26499
rect 14531 26427 14716 26465
rect 14531 26393 14606 26427
rect 14640 26393 14716 26427
rect 14531 26355 14716 26393
rect 14531 26321 14606 26355
rect 14640 26321 14716 26355
rect 14531 26283 14716 26321
rect 14531 26249 14606 26283
rect 14640 26249 14716 26283
rect 14531 26211 14716 26249
rect 14531 26177 14606 26211
rect 14640 26177 14716 26211
rect 14531 26139 14716 26177
rect 14531 26105 14606 26139
rect 14640 26105 14716 26139
rect 14531 26067 14716 26105
rect 14531 26033 14606 26067
rect 14640 26033 14716 26067
rect 14531 25995 14716 26033
rect 14531 25961 14606 25995
rect 14640 25961 14716 25995
rect 14531 25923 14716 25961
rect 14531 25889 14606 25923
rect 14640 25889 14716 25923
rect 14531 25851 14716 25889
rect 14531 25817 14606 25851
rect 14640 25817 14716 25851
rect 14531 25779 14716 25817
rect 14531 25745 14606 25779
rect 14640 25745 14716 25779
rect 14531 25707 14716 25745
rect 14531 25673 14606 25707
rect 14640 25673 14716 25707
rect 14531 25635 14716 25673
rect 14531 25601 14606 25635
rect 14640 25601 14716 25635
rect 14531 25563 14716 25601
rect 14531 25529 14606 25563
rect 14640 25529 14716 25563
rect 14531 25491 14716 25529
rect 14531 25457 14606 25491
rect 14640 25457 14716 25491
rect 14531 25419 14716 25457
rect 14531 25385 14606 25419
rect 14640 25385 14716 25419
rect 14531 25347 14716 25385
rect 14531 25313 14606 25347
rect 14640 25313 14716 25347
rect 14531 25275 14716 25313
rect 14531 25241 14606 25275
rect 14640 25241 14716 25275
rect 14531 25203 14716 25241
rect 14531 25169 14606 25203
rect 14640 25169 14716 25203
rect 14531 25131 14716 25169
rect 14531 25097 14606 25131
rect 14640 25097 14716 25131
rect 14531 25059 14716 25097
rect 14531 25025 14606 25059
rect 14640 25025 14716 25059
rect 14531 24987 14716 25025
rect 14531 24953 14606 24987
rect 14640 24953 14716 24987
rect 14531 24915 14716 24953
rect 14531 24881 14606 24915
rect 14640 24881 14716 24915
rect 14531 24843 14716 24881
rect 14531 24809 14606 24843
rect 14640 24809 14716 24843
rect 14531 24771 14716 24809
rect 14531 24737 14606 24771
rect 14640 24737 14716 24771
rect 14531 24699 14716 24737
rect 14531 24665 14606 24699
rect 14640 24665 14716 24699
rect 14531 24627 14716 24665
rect 14531 24593 14606 24627
rect 14640 24593 14716 24627
rect 14531 24555 14716 24593
rect 14531 24521 14606 24555
rect 14640 24521 14716 24555
rect 14531 24483 14716 24521
rect 14531 24449 14606 24483
rect 14640 24449 14716 24483
rect 14531 24411 14716 24449
rect 14531 24377 14606 24411
rect 14640 24377 14716 24411
rect 14531 24339 14716 24377
rect 14531 24305 14606 24339
rect 14640 24305 14716 24339
rect 14531 24267 14716 24305
rect 14531 24233 14606 24267
rect 14640 24233 14716 24267
rect 14531 24195 14716 24233
rect 14531 24161 14606 24195
rect 14640 24161 14716 24195
rect 14531 24123 14716 24161
rect 14531 24089 14606 24123
rect 14640 24089 14716 24123
rect 14531 24051 14716 24089
rect 14531 24017 14606 24051
rect 14640 24017 14716 24051
rect 14531 23979 14716 24017
rect 14531 23945 14606 23979
rect 14640 23945 14716 23979
rect 14531 23907 14716 23945
rect 14531 23873 14606 23907
rect 14640 23873 14716 23907
rect 14531 23835 14716 23873
rect 14531 23801 14606 23835
rect 14640 23801 14716 23835
rect 14531 23763 14716 23801
rect 14531 23729 14606 23763
rect 14640 23729 14716 23763
rect 14531 23691 14716 23729
rect 14531 23657 14606 23691
rect 14640 23657 14716 23691
rect 14531 23619 14716 23657
rect 14531 23585 14606 23619
rect 14640 23585 14716 23619
rect 14531 23547 14716 23585
rect 14531 23513 14606 23547
rect 14640 23513 14716 23547
rect 14531 23475 14716 23513
rect 14531 23441 14606 23475
rect 14640 23441 14716 23475
rect 14531 23403 14716 23441
rect 14531 23369 14606 23403
rect 14640 23369 14716 23403
rect 14531 23331 14716 23369
rect 14531 23297 14606 23331
rect 14640 23297 14716 23331
rect 14531 23259 14716 23297
rect 14531 23225 14606 23259
rect 14640 23225 14716 23259
rect 14531 23187 14716 23225
rect 14531 23153 14606 23187
rect 14640 23153 14716 23187
rect 14531 23115 14716 23153
rect 14531 23081 14606 23115
rect 14640 23081 14716 23115
rect 14531 23043 14716 23081
rect 14531 23009 14606 23043
rect 14640 23009 14716 23043
rect 14531 22971 14716 23009
rect 14531 22937 14606 22971
rect 14640 22937 14716 22971
rect 14531 22899 14716 22937
rect 14531 22865 14606 22899
rect 14640 22865 14716 22899
rect 14531 22827 14716 22865
rect 14531 22793 14606 22827
rect 14640 22793 14716 22827
rect 14531 22755 14716 22793
rect 14531 22721 14606 22755
rect 14640 22721 14716 22755
rect 14531 22683 14716 22721
rect 14531 22649 14606 22683
rect 14640 22649 14716 22683
rect 14531 22611 14716 22649
rect 14531 22577 14606 22611
rect 14640 22577 14716 22611
rect 14531 22539 14716 22577
rect 14531 22505 14606 22539
rect 14640 22505 14716 22539
rect 14531 22467 14716 22505
rect 14531 22433 14606 22467
rect 14640 22433 14716 22467
rect 14531 22395 14716 22433
rect 14531 22361 14606 22395
rect 14640 22361 14716 22395
rect 14531 22323 14716 22361
rect 14531 22289 14606 22323
rect 14640 22289 14716 22323
rect 14531 22251 14716 22289
rect 14531 22217 14606 22251
rect 14640 22217 14716 22251
rect 14531 22179 14716 22217
rect 14531 22145 14606 22179
rect 14640 22145 14716 22179
rect 14531 22107 14716 22145
rect 14531 22073 14606 22107
rect 14640 22073 14716 22107
rect 14531 22035 14716 22073
rect 14531 22001 14606 22035
rect 14640 22001 14716 22035
rect 14531 21963 14716 22001
rect 14531 21929 14606 21963
rect 14640 21929 14716 21963
rect 14531 21891 14716 21929
rect 14531 21857 14606 21891
rect 14640 21857 14716 21891
rect 14531 21819 14716 21857
rect 14531 21785 14606 21819
rect 14640 21785 14716 21819
rect 14531 21747 14716 21785
rect 14531 21713 14606 21747
rect 14640 21713 14716 21747
rect 14531 21675 14716 21713
rect 14531 21641 14606 21675
rect 14640 21641 14716 21675
rect 14531 21603 14716 21641
rect 14531 21569 14606 21603
rect 14640 21569 14716 21603
rect 14531 21531 14716 21569
rect 14531 21497 14606 21531
rect 14640 21497 14716 21531
rect 14531 21459 14716 21497
rect 14531 21425 14606 21459
rect 14640 21425 14716 21459
rect 14531 21387 14716 21425
rect 14531 21353 14606 21387
rect 14640 21353 14716 21387
rect 14531 21315 14716 21353
rect 14531 21281 14606 21315
rect 14640 21281 14716 21315
rect 14531 21243 14716 21281
rect 14531 21209 14606 21243
rect 14640 21209 14716 21243
rect 14531 21171 14716 21209
rect 14531 21137 14606 21171
rect 14640 21137 14716 21171
rect 14531 21099 14716 21137
rect 14531 21065 14606 21099
rect 14640 21065 14716 21099
rect 14531 21027 14716 21065
rect 14531 20993 14606 21027
rect 14640 20993 14716 21027
rect 14531 20955 14716 20993
rect 14531 20921 14606 20955
rect 14640 20921 14716 20955
rect 14531 20883 14716 20921
rect 14531 20849 14606 20883
rect 14640 20849 14716 20883
rect 14531 20811 14716 20849
rect 14531 20777 14606 20811
rect 14640 20777 14716 20811
rect 14531 20739 14716 20777
rect 14531 20705 14606 20739
rect 14640 20705 14716 20739
rect 14531 20667 14716 20705
rect 14531 20633 14606 20667
rect 14640 20633 14716 20667
rect 14531 20595 14716 20633
rect 14531 20561 14606 20595
rect 14640 20561 14716 20595
rect 14531 20523 14716 20561
rect 14531 20489 14606 20523
rect 14640 20489 14716 20523
rect 14531 20451 14716 20489
rect 14531 20417 14606 20451
rect 14640 20417 14716 20451
rect 14531 20379 14716 20417
rect 14531 20345 14606 20379
rect 14640 20345 14716 20379
rect 14531 20307 14716 20345
rect 14531 20273 14606 20307
rect 14640 20273 14716 20307
rect 14531 20235 14716 20273
rect 14531 20201 14606 20235
rect 14640 20201 14716 20235
rect 14531 20163 14716 20201
rect 14531 20129 14606 20163
rect 14640 20129 14716 20163
rect 14531 20091 14716 20129
rect 14531 20057 14606 20091
rect 14640 20057 14716 20091
rect 14531 20019 14716 20057
rect 14531 19985 14606 20019
rect 14640 19985 14716 20019
rect 14531 19947 14716 19985
rect 14531 19913 14606 19947
rect 14640 19913 14716 19947
rect 14531 19875 14716 19913
rect 14531 19841 14606 19875
rect 14640 19841 14716 19875
rect 14531 19803 14716 19841
rect 14531 19769 14606 19803
rect 14640 19769 14716 19803
rect 14531 19731 14716 19769
rect 14531 19697 14606 19731
rect 14640 19697 14716 19731
rect 14531 19659 14716 19697
rect 14531 19625 14606 19659
rect 14640 19625 14716 19659
rect 14531 19587 14716 19625
rect 14531 19553 14606 19587
rect 14640 19553 14716 19587
rect 14531 19515 14716 19553
rect 14531 19481 14606 19515
rect 14640 19481 14716 19515
rect 14531 19443 14716 19481
rect 14531 19409 14606 19443
rect 14640 19409 14716 19443
rect 14531 19371 14716 19409
rect 14531 19337 14606 19371
rect 14640 19337 14716 19371
rect 14531 19299 14716 19337
rect 14531 19265 14606 19299
rect 14640 19265 14716 19299
rect 14531 19227 14716 19265
rect 14531 19193 14606 19227
rect 14640 19193 14716 19227
rect 14531 19155 14716 19193
rect 14531 19121 14606 19155
rect 14640 19121 14716 19155
rect 14531 19083 14716 19121
rect 14531 19049 14606 19083
rect 14640 19049 14716 19083
rect 14531 19011 14716 19049
rect 14531 18977 14606 19011
rect 14640 18977 14716 19011
rect 14531 18939 14716 18977
rect 14531 18905 14606 18939
rect 14640 18905 14716 18939
rect 14531 18867 14716 18905
rect 14531 18833 14606 18867
rect 14640 18833 14716 18867
rect 14531 18795 14716 18833
rect 14531 18761 14606 18795
rect 14640 18761 14716 18795
rect 14531 18723 14716 18761
rect 14531 18689 14606 18723
rect 14640 18689 14716 18723
rect 14531 18651 14716 18689
rect 14531 18617 14606 18651
rect 14640 18617 14716 18651
rect 14531 18579 14716 18617
rect 14531 18545 14606 18579
rect 14640 18545 14716 18579
rect 14531 18507 14716 18545
rect 14531 18473 14606 18507
rect 14640 18473 14716 18507
rect 14531 18435 14716 18473
rect 14531 18401 14606 18435
rect 14640 18401 14716 18435
rect 14531 18363 14716 18401
rect 14531 18329 14606 18363
rect 14640 18329 14716 18363
rect 14531 18291 14716 18329
rect 14531 18257 14606 18291
rect 14640 18257 14716 18291
rect 14531 18219 14716 18257
rect 14531 18185 14606 18219
rect 14640 18185 14716 18219
rect 14531 18147 14716 18185
rect 14531 18113 14606 18147
rect 14640 18113 14716 18147
rect 14531 18075 14716 18113
rect 14531 18041 14606 18075
rect 14640 18041 14716 18075
rect 14531 18003 14716 18041
rect 14531 17969 14606 18003
rect 14640 17969 14716 18003
rect 14531 17931 14716 17969
rect 14531 17897 14606 17931
rect 14640 17897 14716 17931
rect 14531 17859 14716 17897
rect 14531 17825 14606 17859
rect 14640 17825 14716 17859
rect 14531 17787 14716 17825
rect 14531 17753 14606 17787
rect 14640 17753 14716 17787
rect 14531 17715 14716 17753
rect 14531 17681 14606 17715
rect 14640 17681 14716 17715
rect 14531 17643 14716 17681
rect 14531 17609 14606 17643
rect 14640 17609 14716 17643
rect 14531 17571 14716 17609
rect 14531 17537 14606 17571
rect 14640 17537 14716 17571
rect 14531 17499 14716 17537
rect 14531 17465 14606 17499
rect 14640 17465 14716 17499
rect 14531 17427 14716 17465
rect 14531 17393 14606 17427
rect 14640 17393 14716 17427
rect 14531 17355 14716 17393
rect 14531 17321 14606 17355
rect 14640 17321 14716 17355
rect 14531 17283 14716 17321
rect 14531 17249 14606 17283
rect 14640 17249 14716 17283
rect 14531 17211 14716 17249
rect 14531 17177 14606 17211
rect 14640 17177 14716 17211
rect 14531 17139 14716 17177
rect 14531 17105 14606 17139
rect 14640 17105 14716 17139
rect 14531 17067 14716 17105
rect 14531 17033 14606 17067
rect 14640 17033 14716 17067
rect 14531 16995 14716 17033
rect 14531 16961 14606 16995
rect 14640 16961 14716 16995
rect 14531 16923 14716 16961
rect 14531 16889 14606 16923
rect 14640 16889 14716 16923
rect 14531 16851 14716 16889
rect 14531 16817 14606 16851
rect 14640 16817 14716 16851
rect 14531 16779 14716 16817
rect 14531 16745 14606 16779
rect 14640 16745 14716 16779
rect 14531 16707 14716 16745
rect 14531 16673 14606 16707
rect 14640 16673 14716 16707
rect 14531 16635 14716 16673
rect 14531 16601 14606 16635
rect 14640 16601 14716 16635
rect 14531 16563 14716 16601
rect 14531 16529 14606 16563
rect 14640 16529 14716 16563
rect 14531 16491 14716 16529
rect 14531 16457 14606 16491
rect 14640 16457 14716 16491
rect 14531 16419 14716 16457
rect 14531 16385 14606 16419
rect 14640 16385 14716 16419
rect 14531 16347 14716 16385
rect 14531 16313 14606 16347
rect 14640 16313 14716 16347
rect 14531 16275 14716 16313
rect 14531 16241 14606 16275
rect 14640 16241 14716 16275
rect 14531 16203 14716 16241
rect 14531 16169 14606 16203
rect 14640 16169 14716 16203
rect 14531 16131 14716 16169
rect 14531 16097 14606 16131
rect 14640 16097 14716 16131
rect 14531 16059 14716 16097
rect 14531 16025 14606 16059
rect 14640 16025 14716 16059
rect 14531 15987 14716 16025
rect 14531 15953 14606 15987
rect 14640 15953 14716 15987
rect 14531 15915 14716 15953
rect 14531 15881 14606 15915
rect 14640 15881 14716 15915
rect 14531 15843 14716 15881
rect 14531 15809 14606 15843
rect 14640 15809 14716 15843
rect 14531 15771 14716 15809
rect 14531 15737 14606 15771
rect 14640 15737 14716 15771
rect 14531 15699 14716 15737
rect 14531 15665 14606 15699
rect 14640 15665 14716 15699
rect 14531 15627 14716 15665
rect 14531 15593 14606 15627
rect 14640 15593 14716 15627
rect 14531 15555 14716 15593
rect 14531 15521 14606 15555
rect 14640 15521 14716 15555
rect 14531 15483 14716 15521
rect 14531 15449 14606 15483
rect 14640 15449 14716 15483
rect 14531 15411 14716 15449
rect 14531 15377 14606 15411
rect 14640 15377 14716 15411
rect 14531 15339 14716 15377
rect 14531 15305 14606 15339
rect 14640 15305 14716 15339
rect 14531 15267 14716 15305
rect 14531 15233 14606 15267
rect 14640 15233 14716 15267
rect 14531 15195 14716 15233
rect 14531 15161 14606 15195
rect 14640 15161 14716 15195
rect 14531 15123 14716 15161
rect 14531 15089 14606 15123
rect 14640 15089 14716 15123
rect 14531 15051 14716 15089
rect 14531 15017 14606 15051
rect 14640 15017 14716 15051
rect 14531 14979 14716 15017
rect 14531 14945 14606 14979
rect 14640 14945 14716 14979
rect 14531 14907 14716 14945
rect 14531 14873 14606 14907
rect 14640 14873 14716 14907
rect 237 14804 312 14838
rect 346 14804 422 14838
rect 237 14766 422 14804
rect 237 14732 312 14766
rect 346 14732 422 14766
rect 237 14694 422 14732
rect 237 14660 312 14694
rect 346 14660 422 14694
rect 237 14541 422 14660
rect 850 14787 2088 14856
rect 850 14753 875 14787
rect 909 14753 947 14787
rect 981 14753 1019 14787
rect 1053 14753 1091 14787
rect 1125 14753 1163 14787
rect 1197 14753 1235 14787
rect 1269 14753 1307 14787
rect 1341 14753 1379 14787
rect 1413 14753 1451 14787
rect 1485 14753 1523 14787
rect 1557 14753 1595 14787
rect 1629 14753 1667 14787
rect 1701 14753 1739 14787
rect 1773 14753 1811 14787
rect 1845 14753 1883 14787
rect 1917 14753 1955 14787
rect 1989 14753 2027 14787
rect 2061 14753 2088 14787
rect 850 14744 2088 14753
rect 237 14465 712 14541
rect 237 14431 312 14465
rect 346 14431 602 14465
rect 636 14431 712 14465
rect 237 14356 712 14431
rect 850 14308 900 14744
rect 2040 14308 2088 14744
rect 12850 14787 14088 14856
rect 12850 14753 12875 14787
rect 12909 14753 12947 14787
rect 12981 14753 13019 14787
rect 13053 14753 13091 14787
rect 13125 14753 13163 14787
rect 13197 14753 13235 14787
rect 13269 14753 13307 14787
rect 13341 14753 13379 14787
rect 13413 14753 13451 14787
rect 13485 14753 13523 14787
rect 13557 14753 13595 14787
rect 13629 14753 13667 14787
rect 13701 14753 13739 14787
rect 13773 14753 13811 14787
rect 13845 14753 13883 14787
rect 13917 14753 13955 14787
rect 13989 14753 14027 14787
rect 14061 14753 14088 14787
rect 12850 14744 14088 14753
rect 2240 14465 12697 14541
rect 2240 14431 2303 14465
rect 2337 14431 2375 14465
rect 2409 14431 2447 14465
rect 2481 14431 2519 14465
rect 2553 14431 2591 14465
rect 2625 14431 2663 14465
rect 2697 14431 2735 14465
rect 2769 14431 2807 14465
rect 2841 14431 2879 14465
rect 2913 14431 2951 14465
rect 2985 14431 3023 14465
rect 3057 14431 3095 14465
rect 3129 14431 3167 14465
rect 3201 14431 3239 14465
rect 3273 14431 3311 14465
rect 3345 14431 3383 14465
rect 3417 14431 3455 14465
rect 3489 14431 3527 14465
rect 3561 14431 3599 14465
rect 3633 14431 3671 14465
rect 3705 14431 3743 14465
rect 3777 14431 3815 14465
rect 3849 14431 3887 14465
rect 3921 14431 3959 14465
rect 3993 14431 4031 14465
rect 4065 14431 4103 14465
rect 4137 14431 4175 14465
rect 4209 14431 4247 14465
rect 4281 14431 4319 14465
rect 4353 14431 4391 14465
rect 4425 14431 4463 14465
rect 4497 14431 4535 14465
rect 4569 14431 4607 14465
rect 4641 14431 4679 14465
rect 4713 14431 4751 14465
rect 4785 14431 4823 14465
rect 4857 14431 4895 14465
rect 4929 14431 4967 14465
rect 5001 14431 5039 14465
rect 5073 14431 5111 14465
rect 5145 14431 5183 14465
rect 5217 14431 5255 14465
rect 5289 14431 5327 14465
rect 5361 14431 5399 14465
rect 5433 14431 5471 14465
rect 5505 14431 5543 14465
rect 5577 14431 5615 14465
rect 5649 14431 5687 14465
rect 5721 14431 5759 14465
rect 5793 14431 5831 14465
rect 5865 14431 5903 14465
rect 5937 14431 5975 14465
rect 6009 14431 6047 14465
rect 6081 14431 6119 14465
rect 6153 14431 6191 14465
rect 6225 14431 6263 14465
rect 6297 14431 6335 14465
rect 6369 14431 6407 14465
rect 6441 14431 6479 14465
rect 6513 14431 6551 14465
rect 6585 14431 6623 14465
rect 6657 14431 6695 14465
rect 6729 14431 6767 14465
rect 6801 14431 6839 14465
rect 6873 14431 6911 14465
rect 6945 14431 6983 14465
rect 7017 14431 7055 14465
rect 7089 14431 7127 14465
rect 7161 14431 7199 14465
rect 7233 14431 7271 14465
rect 7305 14431 7343 14465
rect 7377 14431 7415 14465
rect 7449 14431 7487 14465
rect 7521 14431 7559 14465
rect 7593 14431 7631 14465
rect 7665 14431 7703 14465
rect 7737 14431 7775 14465
rect 7809 14431 7847 14465
rect 7881 14431 7919 14465
rect 7953 14431 7991 14465
rect 8025 14431 8063 14465
rect 8097 14431 8135 14465
rect 8169 14431 8207 14465
rect 8241 14431 8279 14465
rect 8313 14431 8351 14465
rect 8385 14431 8423 14465
rect 8457 14431 8495 14465
rect 8529 14431 8567 14465
rect 8601 14431 8639 14465
rect 8673 14431 8711 14465
rect 8745 14431 8783 14465
rect 8817 14431 8855 14465
rect 8889 14431 8927 14465
rect 8961 14431 8999 14465
rect 9033 14431 9071 14465
rect 9105 14431 9143 14465
rect 9177 14431 9215 14465
rect 9249 14431 9287 14465
rect 9321 14431 9359 14465
rect 9393 14431 9431 14465
rect 9465 14431 9503 14465
rect 9537 14431 9575 14465
rect 9609 14431 9647 14465
rect 9681 14431 9719 14465
rect 9753 14431 9791 14465
rect 9825 14431 9863 14465
rect 9897 14431 9935 14465
rect 9969 14431 10007 14465
rect 10041 14431 10079 14465
rect 10113 14431 10151 14465
rect 10185 14431 10223 14465
rect 10257 14431 10295 14465
rect 10329 14431 10367 14465
rect 10401 14431 10439 14465
rect 10473 14431 10511 14465
rect 10545 14431 10583 14465
rect 10617 14431 10655 14465
rect 10689 14431 10727 14465
rect 10761 14431 10799 14465
rect 10833 14431 10871 14465
rect 10905 14431 10943 14465
rect 10977 14431 11015 14465
rect 11049 14431 11087 14465
rect 11121 14431 11159 14465
rect 11193 14431 11231 14465
rect 11265 14431 11303 14465
rect 11337 14431 11375 14465
rect 11409 14431 11447 14465
rect 11481 14431 11519 14465
rect 11553 14431 11591 14465
rect 11625 14431 11663 14465
rect 11697 14431 11735 14465
rect 11769 14431 11807 14465
rect 11841 14431 11879 14465
rect 11913 14431 11951 14465
rect 11985 14431 12023 14465
rect 12057 14431 12095 14465
rect 12129 14431 12167 14465
rect 12201 14431 12239 14465
rect 12273 14431 12311 14465
rect 12345 14431 12383 14465
rect 12417 14431 12455 14465
rect 12489 14431 12527 14465
rect 12561 14431 12599 14465
rect 12633 14431 12697 14465
rect 2240 14356 12697 14431
rect 850 14265 2088 14308
rect 12850 14308 12900 14744
rect 14040 14308 14088 14744
rect 14531 14835 14716 14873
rect 14531 14801 14606 14835
rect 14640 14801 14716 14835
rect 14531 14763 14716 14801
rect 14531 14729 14606 14763
rect 14640 14729 14716 14763
rect 14531 14691 14716 14729
rect 14531 14657 14606 14691
rect 14640 14657 14716 14691
rect 14531 14541 14716 14657
rect 14224 14465 14716 14541
rect 14224 14431 14306 14465
rect 14340 14431 14606 14465
rect 14640 14431 14716 14465
rect 14224 14356 14716 14431
rect 12850 14265 14088 14308
<< via1 >>
rect 949 36511 2153 37224
rect 12813 36511 14017 37221
rect 949 36477 980 36511
rect 980 36477 1014 36511
rect 1014 36477 1052 36511
rect 1052 36477 1086 36511
rect 1086 36477 1124 36511
rect 1124 36477 1158 36511
rect 1158 36477 1196 36511
rect 1196 36477 1230 36511
rect 1230 36477 1268 36511
rect 1268 36477 1302 36511
rect 1302 36477 1340 36511
rect 1340 36477 1374 36511
rect 1374 36477 1412 36511
rect 1412 36477 1446 36511
rect 1446 36477 1484 36511
rect 1484 36477 1518 36511
rect 1518 36477 1556 36511
rect 1556 36477 1590 36511
rect 1590 36477 1628 36511
rect 1628 36477 1662 36511
rect 1662 36477 1700 36511
rect 1700 36477 1734 36511
rect 1734 36477 1772 36511
rect 1772 36477 1806 36511
rect 1806 36477 1844 36511
rect 1844 36477 1878 36511
rect 1878 36477 1916 36511
rect 1916 36477 1950 36511
rect 1950 36477 1988 36511
rect 1988 36477 2022 36511
rect 2022 36477 2060 36511
rect 2060 36477 2094 36511
rect 2094 36477 2132 36511
rect 2132 36477 2153 36511
rect 12813 36477 12822 36511
rect 12822 36477 12860 36511
rect 12860 36477 12894 36511
rect 12894 36477 12932 36511
rect 12932 36477 12966 36511
rect 12966 36477 13004 36511
rect 13004 36477 13038 36511
rect 13038 36477 13076 36511
rect 13076 36477 13110 36511
rect 13110 36477 13148 36511
rect 13148 36477 13182 36511
rect 13182 36477 13220 36511
rect 13220 36477 13254 36511
rect 13254 36477 13292 36511
rect 13292 36477 13326 36511
rect 13326 36477 13364 36511
rect 13364 36477 13398 36511
rect 13398 36477 13436 36511
rect 13436 36477 13470 36511
rect 13470 36477 13508 36511
rect 13508 36477 13542 36511
rect 13542 36477 13580 36511
rect 13580 36477 13614 36511
rect 13614 36477 13652 36511
rect 13652 36477 13686 36511
rect 13686 36477 13724 36511
rect 13724 36477 13758 36511
rect 13758 36477 13796 36511
rect 13796 36477 13830 36511
rect 13830 36477 13868 36511
rect 13868 36477 13902 36511
rect 13902 36477 13940 36511
rect 13940 36477 13974 36511
rect 13974 36477 14012 36511
rect 14012 36477 14017 36511
rect 949 36468 2153 36477
rect 12813 36465 14017 36477
rect 4936 29420 7228 30240
rect 7737 29420 10029 30240
rect 4931 28277 7223 28348
rect 7742 28277 10034 28348
rect 4931 28243 4963 28277
rect 4963 28243 4997 28277
rect 4997 28243 5035 28277
rect 5035 28243 5069 28277
rect 5069 28243 5107 28277
rect 5107 28243 5141 28277
rect 5141 28243 5179 28277
rect 5179 28243 5213 28277
rect 5213 28243 5251 28277
rect 5251 28243 5285 28277
rect 5285 28243 5323 28277
rect 5323 28243 5357 28277
rect 5357 28243 5395 28277
rect 5395 28243 5429 28277
rect 5429 28243 5467 28277
rect 5467 28243 5501 28277
rect 5501 28243 5539 28277
rect 5539 28243 5573 28277
rect 5573 28243 5611 28277
rect 5611 28243 5645 28277
rect 5645 28243 5683 28277
rect 5683 28243 5717 28277
rect 5717 28243 5755 28277
rect 5755 28243 5789 28277
rect 5789 28243 5827 28277
rect 5827 28243 5861 28277
rect 5861 28243 5899 28277
rect 5899 28243 5933 28277
rect 5933 28243 5971 28277
rect 5971 28243 6005 28277
rect 6005 28243 6043 28277
rect 6043 28243 6077 28277
rect 6077 28243 6115 28277
rect 6115 28243 6149 28277
rect 6149 28243 6187 28277
rect 6187 28243 6221 28277
rect 6221 28243 6259 28277
rect 6259 28243 6293 28277
rect 6293 28243 6331 28277
rect 6331 28243 6365 28277
rect 6365 28243 6403 28277
rect 6403 28243 6437 28277
rect 6437 28243 6475 28277
rect 6475 28243 6509 28277
rect 6509 28243 6547 28277
rect 6547 28243 6581 28277
rect 6581 28243 6619 28277
rect 6619 28243 6653 28277
rect 6653 28243 6691 28277
rect 6691 28243 6725 28277
rect 6725 28243 6763 28277
rect 6763 28243 6797 28277
rect 6797 28243 6835 28277
rect 6835 28243 6869 28277
rect 6869 28243 6907 28277
rect 6907 28243 6941 28277
rect 6941 28243 6979 28277
rect 6979 28243 7013 28277
rect 7013 28243 7051 28277
rect 7051 28243 7085 28277
rect 7085 28243 7123 28277
rect 7123 28243 7157 28277
rect 7157 28243 7195 28277
rect 7195 28243 7223 28277
rect 7742 28243 7771 28277
rect 7771 28243 7805 28277
rect 7805 28243 7843 28277
rect 7843 28243 7877 28277
rect 7877 28243 7915 28277
rect 7915 28243 7949 28277
rect 7949 28243 7987 28277
rect 7987 28243 8021 28277
rect 8021 28243 8059 28277
rect 8059 28243 8093 28277
rect 8093 28243 8131 28277
rect 8131 28243 8165 28277
rect 8165 28243 8203 28277
rect 8203 28243 8237 28277
rect 8237 28243 8275 28277
rect 8275 28243 8309 28277
rect 8309 28243 8347 28277
rect 8347 28243 8381 28277
rect 8381 28243 8419 28277
rect 8419 28243 8453 28277
rect 8453 28243 8491 28277
rect 8491 28243 8525 28277
rect 8525 28243 8563 28277
rect 8563 28243 8597 28277
rect 8597 28243 8635 28277
rect 8635 28243 8669 28277
rect 8669 28243 8707 28277
rect 8707 28243 8741 28277
rect 8741 28243 8779 28277
rect 8779 28243 8813 28277
rect 8813 28243 8851 28277
rect 8851 28243 8885 28277
rect 8885 28243 8923 28277
rect 8923 28243 8957 28277
rect 8957 28243 8995 28277
rect 8995 28243 9029 28277
rect 9029 28243 9067 28277
rect 9067 28243 9101 28277
rect 9101 28243 9139 28277
rect 9139 28243 9173 28277
rect 9173 28243 9211 28277
rect 9211 28243 9245 28277
rect 9245 28243 9283 28277
rect 9283 28243 9317 28277
rect 9317 28243 9355 28277
rect 9355 28243 9389 28277
rect 9389 28243 9427 28277
rect 9427 28243 9461 28277
rect 9461 28243 9499 28277
rect 9499 28243 9533 28277
rect 9533 28243 9571 28277
rect 9571 28243 9605 28277
rect 9605 28243 9643 28277
rect 9643 28243 9677 28277
rect 9677 28243 9715 28277
rect 9715 28243 9749 28277
rect 9749 28243 9787 28277
rect 9787 28243 9821 28277
rect 9821 28243 9859 28277
rect 9859 28243 9893 28277
rect 9893 28243 9931 28277
rect 9931 28243 9965 28277
rect 9965 28243 10003 28277
rect 10003 28243 10034 28277
rect 4931 28232 7223 28243
rect 7742 28232 10034 28243
rect 2501 28032 4473 28035
rect 10492 28032 12464 28035
rect 2501 27926 2515 28032
rect 2515 27926 4473 28032
rect 10492 27926 12464 28032
rect 2501 27919 4473 27926
rect 10492 27919 12464 27926
rect 4931 27683 7223 27732
rect 7742 27683 10034 27732
rect 4931 27616 7223 27683
rect 7742 27616 10034 27683
rect 4925 25922 7217 26038
rect 7749 25922 10041 26038
rect 2538 25760 4446 25772
rect 10520 25760 12428 25772
rect 2538 25656 4446 25760
rect 10520 25656 12428 25760
rect 4925 25505 4951 25506
rect 4951 25505 4985 25506
rect 4985 25505 5023 25506
rect 5023 25505 5057 25506
rect 5057 25505 5095 25506
rect 5095 25505 5129 25506
rect 5129 25505 5167 25506
rect 5167 25505 5201 25506
rect 5201 25505 5239 25506
rect 5239 25505 5273 25506
rect 5273 25505 5311 25506
rect 5311 25505 5345 25506
rect 5345 25505 5383 25506
rect 5383 25505 5417 25506
rect 5417 25505 5455 25506
rect 5455 25505 5489 25506
rect 5489 25505 5527 25506
rect 5527 25505 5561 25506
rect 5561 25505 5599 25506
rect 5599 25505 5633 25506
rect 5633 25505 5671 25506
rect 5671 25505 5705 25506
rect 5705 25505 5743 25506
rect 5743 25505 5777 25506
rect 5777 25505 5815 25506
rect 5815 25505 5849 25506
rect 5849 25505 5887 25506
rect 5887 25505 5921 25506
rect 5921 25505 5959 25506
rect 5959 25505 5993 25506
rect 5993 25505 6031 25506
rect 6031 25505 6065 25506
rect 6065 25505 6103 25506
rect 6103 25505 6137 25506
rect 6137 25505 6175 25506
rect 6175 25505 6209 25506
rect 6209 25505 6247 25506
rect 6247 25505 6281 25506
rect 6281 25505 6319 25506
rect 6319 25505 6353 25506
rect 6353 25505 6391 25506
rect 6391 25505 6425 25506
rect 6425 25505 6463 25506
rect 6463 25505 6497 25506
rect 6497 25505 6535 25506
rect 6535 25505 6569 25506
rect 6569 25505 6607 25506
rect 6607 25505 6641 25506
rect 6641 25505 6679 25506
rect 6679 25505 6713 25506
rect 6713 25505 6751 25506
rect 6751 25505 6785 25506
rect 6785 25505 6823 25506
rect 6823 25505 6857 25506
rect 6857 25505 6895 25506
rect 6895 25505 6929 25506
rect 6929 25505 6967 25506
rect 6967 25505 7001 25506
rect 7001 25505 7039 25506
rect 7039 25505 7073 25506
rect 7073 25505 7111 25506
rect 7111 25505 7145 25506
rect 7145 25505 7183 25506
rect 7183 25505 7217 25506
rect 7749 25505 7759 25506
rect 7759 25505 7793 25506
rect 7793 25505 7831 25506
rect 7831 25505 7865 25506
rect 7865 25505 7903 25506
rect 7903 25505 7937 25506
rect 7937 25505 7975 25506
rect 7975 25505 8009 25506
rect 8009 25505 8047 25506
rect 8047 25505 8081 25506
rect 8081 25505 8119 25506
rect 8119 25505 8153 25506
rect 8153 25505 8191 25506
rect 8191 25505 8225 25506
rect 8225 25505 8263 25506
rect 8263 25505 8297 25506
rect 8297 25505 8335 25506
rect 8335 25505 8369 25506
rect 8369 25505 8407 25506
rect 8407 25505 8441 25506
rect 8441 25505 8479 25506
rect 8479 25505 8513 25506
rect 8513 25505 8551 25506
rect 8551 25505 8585 25506
rect 8585 25505 8623 25506
rect 8623 25505 8657 25506
rect 8657 25505 8695 25506
rect 8695 25505 8729 25506
rect 8729 25505 8767 25506
rect 8767 25505 8801 25506
rect 8801 25505 8839 25506
rect 8839 25505 8873 25506
rect 8873 25505 8911 25506
rect 8911 25505 8945 25506
rect 8945 25505 8983 25506
rect 8983 25505 9017 25506
rect 9017 25505 9055 25506
rect 9055 25505 9089 25506
rect 9089 25505 9127 25506
rect 9127 25505 9161 25506
rect 9161 25505 9199 25506
rect 9199 25505 9233 25506
rect 9233 25505 9271 25506
rect 9271 25505 9305 25506
rect 9305 25505 9343 25506
rect 9343 25505 9377 25506
rect 9377 25505 9415 25506
rect 9415 25505 9449 25506
rect 9449 25505 9487 25506
rect 9487 25505 9521 25506
rect 9521 25505 9559 25506
rect 9559 25505 9593 25506
rect 9593 25505 9631 25506
rect 9631 25505 9665 25506
rect 9665 25505 9703 25506
rect 9703 25505 9737 25506
rect 9737 25505 9775 25506
rect 9775 25505 9809 25506
rect 9809 25505 9847 25506
rect 9847 25505 9881 25506
rect 9881 25505 9919 25506
rect 9919 25505 9953 25506
rect 9953 25505 9991 25506
rect 9991 25505 10025 25506
rect 10025 25505 10041 25506
rect 4925 25390 7217 25505
rect 7749 25390 10041 25505
rect 4937 23682 7229 24502
rect 7736 23682 10028 24502
rect 900 14308 2040 14744
rect 12900 14308 14040 14744
<< metal2 >>
tri 4883 39335 4983 39435 se
rect 4983 39335 7183 39435
tri 7183 39335 7283 39435 sw
rect 4883 39226 7283 39335
rect 877 37224 2226 37271
rect 877 36468 949 37224
rect 2153 36468 2226 37224
rect 877 36421 2226 36468
rect 4883 35330 4971 39226
rect 7187 35330 7283 39226
rect 4883 30240 7283 35330
rect 4883 29420 4936 30240
rect 7228 29420 7283 30240
tri 293 28988 493 29188 se
rect 493 28988 4283 29188
tri 4283 28988 4483 29188 sw
rect 293 28872 4483 28988
rect 293 24816 458 28872
rect 2434 28035 4483 28872
rect 2434 27919 2501 28035
rect 4473 27919 4483 28035
rect 2434 25772 4483 27919
rect 4883 28348 7283 29420
rect 4883 28232 4931 28348
rect 7223 28232 7283 28348
rect 4883 27732 7283 28232
rect 4883 27616 4931 27732
rect 7223 27616 7283 27732
rect 4883 27330 7283 27616
tri 4883 27130 5083 27330 ne
rect 5083 27130 7083 27330
tri 7083 27130 7283 27330 nw
tri 7683 39335 7783 39435 se
rect 7783 39335 9983 39435
tri 9983 39335 10083 39435 sw
rect 7683 39226 10083 39335
rect 7683 35330 7771 39226
rect 9987 35330 10083 39226
rect 12744 37221 14093 37275
rect 12744 36465 12813 37221
rect 14017 36465 14093 37221
rect 12744 36425 14093 36465
rect 7683 30240 10083 35330
rect 7683 29420 7737 30240
rect 10029 29420 10083 30240
rect 7683 28348 10083 29420
rect 7683 28232 7742 28348
rect 10034 28232 10083 28348
rect 7683 27732 10083 28232
rect 7683 27616 7742 27732
rect 10034 27616 10083 27732
rect 7683 27330 10083 27616
tri 7683 27130 7883 27330 ne
rect 7883 27130 9883 27330
tri 9883 27130 10083 27330 nw
tri 10483 28988 10683 29188 se
rect 10683 28988 14423 29188
tri 14423 28988 14623 29188 sw
rect 10483 28920 14623 28988
rect 10483 28035 12447 28920
rect 10483 27919 10492 28035
rect 2434 25656 2538 25772
rect 4446 25656 4483 25772
rect 2434 24816 4483 25656
rect 293 24529 4483 24816
tri 293 24329 493 24529 ne
rect 493 24329 4283 24529
tri 4283 24329 4483 24529 nw
tri 4883 26291 5083 26491 se
rect 5083 26291 7083 26491
tri 7083 26291 7283 26491 sw
rect 4883 26038 7283 26291
rect 4883 25922 4925 26038
rect 7217 25922 7283 26038
rect 4883 25506 7283 25922
rect 4883 25390 4925 25506
rect 7217 25390 7283 25506
rect 4883 24502 7283 25390
rect 4883 23682 4937 24502
rect 7229 23682 7283 24502
tri 2883 19377 4883 21377 se
rect 4883 19377 7283 23682
rect 2883 18944 5283 19377
rect 2883 17288 2934 18944
rect 5230 17288 5283 18944
tri 5283 17377 7283 19377 nw
tri 7683 26291 7883 26491 se
rect 7883 26291 9883 26491
tri 9883 26291 10083 26491 sw
rect 7683 26038 10083 26291
rect 7683 25922 7749 26038
rect 10041 25922 10083 26038
rect 7683 25506 10083 25922
rect 7683 25390 7749 25506
rect 10041 25390 10083 25506
rect 7683 24502 10083 25390
rect 7683 23682 7736 24502
rect 10028 23682 10083 24502
rect 10483 25772 12447 27919
rect 10483 25656 10520 25772
rect 12428 25656 12447 25772
rect 10483 24864 12447 25656
rect 14423 24864 14623 28920
rect 10483 24529 14623 24864
tri 10483 24329 10683 24529 ne
rect 10683 24329 14423 24529
tri 14423 24329 14623 24529 nw
rect 7683 19343 10083 23682
tri 10083 19343 12083 21343 sw
tri 7683 17343 9683 19343 ne
rect 9683 18944 12083 19343
rect 2883 17227 5283 17288
rect 2883 17099 3095 17227
tri 2883 16999 2983 17099 ne
rect 2983 17091 3095 17099
rect 5231 17091 5283 17227
rect 2983 17069 5283 17091
rect 2983 16999 5213 17069
tri 5213 16999 5283 17069 nw
rect 9683 17288 9734 18944
rect 12030 17288 12083 18944
rect 9683 17227 12083 17288
rect 9683 17091 9731 17227
rect 11867 17099 12083 17227
rect 11867 17091 11983 17099
rect 9683 17069 11983 17091
tri 9683 16999 9753 17069 ne
rect 9753 16999 11983 17069
tri 11983 16999 12083 17099 nw
rect 850 14744 2088 14785
rect 850 14308 900 14744
rect 2040 14308 2088 14744
rect 850 14265 2088 14308
rect 12850 14744 14088 14785
rect 12850 14308 12900 14744
rect 14040 14308 14088 14744
rect 12850 14265 14088 14308
<< via2 >>
rect 963 36498 2139 37194
rect 4971 35330 7187 39226
rect 458 24816 2434 28872
rect 7771 35330 9987 39226
rect 12827 36495 14003 37191
rect 12447 28035 14423 28920
rect 12447 27919 12464 28035
rect 12464 27919 14423 28035
rect 2934 17288 5230 18944
rect 12447 24864 14423 27919
rect 3095 17091 5231 17227
rect 9734 17288 12030 18944
rect 9731 17091 11867 17227
<< metal3 >>
tri 4797 39535 5197 39935 se
rect 5197 39870 9778 39935
rect 5197 39566 5259 39870
rect 9723 39566 9778 39870
rect 5197 39535 9778 39566
tri 9778 39535 10178 39935 sw
rect 4797 39468 10178 39535
rect 877 37198 2226 37271
rect 877 36494 959 37198
rect 2143 36494 2226 37198
rect 877 36421 2226 36494
rect 4797 35324 4967 39468
rect 9991 35324 10178 39468
rect 12744 37195 14093 37275
rect 12744 36491 12823 37195
rect 14007 36491 14093 37195
rect 12744 36425 14093 36491
rect 4797 35279 10178 35324
tri 4797 35179 4897 35279 ne
rect 4897 35179 10078 35279
tri 10078 35179 10178 35279 nw
tri 237 33734 1147 34644 se
rect 1147 34588 3092 34644
rect 1147 34124 2331 34588
rect 3035 34124 3092 34588
rect 1147 33861 3092 34124
rect 1147 33734 2692 33861
rect 237 32974 2692 33734
tri 2692 33461 3092 33861 nw
rect 11892 34587 13827 34644
rect 11892 34123 11961 34587
rect 12665 34123 13827 34587
rect 11892 33861 13827 34123
tri 11892 33461 12292 33861 ne
rect 12292 33755 13827 33861
tri 13827 33755 14716 34644 sw
rect 237 28872 1035 32974
rect 1419 28872 2692 32974
rect 237 24816 458 28872
rect 2434 24816 2692 28872
rect 237 21230 1035 24816
rect 1419 21230 2692 24816
rect 237 20451 2692 21230
tri 237 19541 1147 20451 ne
rect 1147 20080 2692 20451
rect 12292 32866 14716 33755
rect 12292 28920 13581 32866
rect 13965 28920 14716 32866
rect 12292 24864 12447 28920
rect 14423 24864 14716 28920
rect 12292 21122 13581 24864
rect 13965 21122 14716 24864
rect 12292 20461 14716 21122
tri 2692 20080 2904 20292 sw
tri 12100 20080 12292 20272 se
rect 12292 20080 13796 20461
rect 1147 20040 13796 20080
rect 1147 19576 2308 20040
rect 12692 19576 13796 20040
rect 1147 19541 13796 19576
tri 13796 19541 14716 20461 nw
tri 2834 19009 3034 19209 se
rect 3034 19009 5372 19209
rect 2834 18944 5372 19009
rect 2834 18908 2934 18944
rect 5230 18908 5372 18944
rect 2834 17324 2930 18908
rect 5234 17324 5372 18908
rect 2834 17288 2934 17324
rect 5230 17288 5372 17324
rect 2834 17243 5372 17288
tri 2834 17043 3034 17243 ne
rect 3034 17231 5372 17243
rect 3034 17087 3091 17231
rect 5235 17087 5372 17231
rect 3034 17043 5372 17087
rect 9588 19009 11927 19209
tri 11927 19009 12127 19209 sw
rect 9588 18944 12127 19009
rect 9588 18908 9734 18944
rect 12030 18908 12127 18944
rect 9588 17324 9730 18908
rect 12034 17324 12127 18908
rect 9588 17288 9734 17324
rect 12030 17288 12127 17324
rect 9588 17243 12127 17288
rect 9588 17231 11927 17243
rect 9588 17087 9727 17231
rect 11871 17087 11927 17231
rect 9588 17043 11927 17087
tri 11927 17043 12127 17243 nw
rect 850 14718 2088 14785
rect 850 14334 918 14718
rect 2022 14334 2088 14718
rect 850 14265 2088 14334
rect 12850 14718 14088 14785
rect 12850 14334 12918 14718
rect 14022 14334 14088 14718
rect 12850 14265 14088 14334
<< via3 >>
rect 5259 39566 9723 39870
rect 959 37194 2143 37198
rect 959 36498 963 37194
rect 963 36498 2139 37194
rect 2139 36498 2143 37194
rect 959 36494 2143 36498
rect 4967 39226 9991 39468
rect 4967 35330 4971 39226
rect 4971 35330 7187 39226
rect 7187 35330 7771 39226
rect 7771 35330 9987 39226
rect 9987 35330 9991 39226
rect 4967 35324 9991 35330
rect 12823 37191 14007 37195
rect 12823 36495 12827 37191
rect 12827 36495 14003 37191
rect 14003 36495 14007 37191
rect 12823 36491 14007 36495
rect 2331 34124 3035 34588
rect 11961 34123 12665 34587
rect 1035 28872 1419 32974
rect 1035 24816 1419 28872
rect 1035 21230 1419 24816
rect 13581 28920 13965 32866
rect 13581 24864 13965 28920
rect 13581 21122 13965 24864
rect 2308 19576 12692 20040
rect 2930 17324 2934 18908
rect 2934 17324 5230 18908
rect 5230 17324 5234 18908
rect 3091 17227 5235 17231
rect 3091 17091 3095 17227
rect 3095 17091 5231 17227
rect 5231 17091 5235 17227
rect 3091 17087 5235 17091
rect 9730 17324 9734 18908
rect 9734 17324 12030 18908
rect 12030 17324 12034 18908
rect 9727 17227 11871 17231
rect 9727 17091 9731 17227
rect 9731 17091 11867 17227
rect 11867 17091 11871 17227
rect 9727 17087 11871 17091
rect 918 14334 2022 14718
rect 12918 14334 14022 14718
<< metal4 >>
rect 0 39965 15000 40000
rect 0 39729 241 39965
rect 477 39729 568 39965
rect 804 39729 895 39965
rect 1131 39729 1222 39965
rect 1458 39729 1549 39965
rect 1785 39729 1876 39965
rect 2112 39729 2203 39965
rect 2439 39729 2530 39965
rect 2766 39729 2857 39965
rect 3093 39729 3184 39965
rect 3420 39729 3511 39965
rect 3747 39729 3838 39965
rect 4074 39729 4165 39965
rect 4401 39729 4492 39965
rect 4728 39729 4819 39965
rect 5055 39729 5146 39965
rect 5382 39870 5473 39965
rect 5709 39870 5800 39965
rect 6036 39870 6127 39965
rect 6363 39870 6454 39965
rect 6690 39870 6781 39965
rect 7017 39870 7108 39965
rect 7344 39870 7435 39965
rect 7671 39870 7762 39965
rect 7998 39870 8089 39965
rect 8325 39870 8415 39965
rect 8651 39870 8741 39965
rect 8977 39870 9067 39965
rect 9303 39870 9393 39965
rect 9629 39870 9719 39965
rect 9955 39729 10045 39965
rect 10281 39729 10371 39965
rect 10607 39729 10697 39965
rect 10933 39729 11023 39965
rect 11259 39729 11349 39965
rect 11585 39729 11675 39965
rect 11911 39729 12001 39965
rect 12237 39729 12327 39965
rect 12563 39729 12653 39965
rect 12889 39729 12979 39965
rect 13215 39729 13305 39965
rect 13541 39729 13631 39965
rect 13867 39729 13957 39965
rect 14193 39729 14283 39965
rect 14519 39729 14609 39965
rect 14845 39729 15000 39965
rect 0 39641 5259 39729
rect 9723 39641 15000 39729
rect 0 39405 241 39641
rect 477 39405 568 39641
rect 804 39405 895 39641
rect 1131 39405 1222 39641
rect 1458 39405 1549 39641
rect 1785 39405 1876 39641
rect 2112 39405 2203 39641
rect 2439 39405 2530 39641
rect 2766 39405 2857 39641
rect 3093 39405 3184 39641
rect 3420 39405 3511 39641
rect 3747 39405 3838 39641
rect 4074 39405 4165 39641
rect 4401 39405 4492 39641
rect 4728 39405 4819 39641
rect 5055 39468 5146 39641
rect 5382 39468 5473 39566
rect 5709 39468 5800 39566
rect 6036 39468 6127 39566
rect 6363 39468 6454 39566
rect 6690 39468 6781 39566
rect 7017 39468 7108 39566
rect 7344 39468 7435 39566
rect 7671 39468 7762 39566
rect 7998 39468 8089 39566
rect 8325 39468 8415 39566
rect 8651 39468 8741 39566
rect 8977 39468 9067 39566
rect 9303 39468 9393 39566
rect 9629 39468 9719 39566
rect 9955 39468 10045 39641
rect 9991 39405 10045 39468
rect 10281 39405 10371 39641
rect 10607 39405 10697 39641
rect 10933 39405 11023 39641
rect 11259 39405 11349 39641
rect 11585 39405 11675 39641
rect 11911 39405 12001 39641
rect 12237 39405 12327 39641
rect 12563 39405 12653 39641
rect 12889 39405 12979 39641
rect 13215 39405 13305 39641
rect 13541 39405 13631 39641
rect 13867 39405 13957 39641
rect 14193 39405 14283 39641
rect 14519 39405 14609 39641
rect 14845 39405 15000 39641
rect 0 39317 4967 39405
rect 9991 39317 15000 39405
rect 0 39081 241 39317
rect 477 39081 568 39317
rect 804 39081 895 39317
rect 1131 39081 1222 39317
rect 1458 39081 1549 39317
rect 1785 39081 1876 39317
rect 2112 39081 2203 39317
rect 2439 39081 2530 39317
rect 2766 39081 2857 39317
rect 3093 39081 3184 39317
rect 3420 39081 3511 39317
rect 3747 39081 3838 39317
rect 4074 39081 4165 39317
rect 4401 39081 4492 39317
rect 4728 39081 4819 39317
rect 9991 39081 10045 39317
rect 10281 39081 10371 39317
rect 10607 39081 10697 39317
rect 10933 39081 11023 39317
rect 11259 39081 11349 39317
rect 11585 39081 11675 39317
rect 11911 39081 12001 39317
rect 12237 39081 12327 39317
rect 12563 39081 12653 39317
rect 12889 39081 12979 39317
rect 13215 39081 13305 39317
rect 13541 39081 13631 39317
rect 13867 39081 13957 39317
rect 14193 39081 14283 39317
rect 14519 39081 14609 39317
rect 14845 39081 15000 39317
rect 0 38993 4967 39081
rect 9991 38993 15000 39081
rect 0 38757 241 38993
rect 477 38757 568 38993
rect 804 38757 895 38993
rect 1131 38757 1222 38993
rect 1458 38757 1549 38993
rect 1785 38757 1876 38993
rect 2112 38757 2203 38993
rect 2439 38757 2530 38993
rect 2766 38757 2857 38993
rect 3093 38757 3184 38993
rect 3420 38757 3511 38993
rect 3747 38757 3838 38993
rect 4074 38757 4165 38993
rect 4401 38757 4492 38993
rect 4728 38757 4819 38993
rect 9991 38757 10045 38993
rect 10281 38757 10371 38993
rect 10607 38757 10697 38993
rect 10933 38757 11023 38993
rect 11259 38757 11349 38993
rect 11585 38757 11675 38993
rect 11911 38757 12001 38993
rect 12237 38757 12327 38993
rect 12563 38757 12653 38993
rect 12889 38757 12979 38993
rect 13215 38757 13305 38993
rect 13541 38757 13631 38993
rect 13867 38757 13957 38993
rect 14193 38757 14283 38993
rect 14519 38757 14609 38993
rect 14845 38757 15000 38993
rect 0 38669 4967 38757
rect 9991 38669 15000 38757
rect 0 38433 241 38669
rect 477 38433 568 38669
rect 804 38433 895 38669
rect 1131 38433 1222 38669
rect 1458 38433 1549 38669
rect 1785 38433 1876 38669
rect 2112 38433 2203 38669
rect 2439 38433 2530 38669
rect 2766 38433 2857 38669
rect 3093 38433 3184 38669
rect 3420 38433 3511 38669
rect 3747 38433 3838 38669
rect 4074 38433 4165 38669
rect 4401 38433 4492 38669
rect 4728 38433 4819 38669
rect 9991 38433 10045 38669
rect 10281 38433 10371 38669
rect 10607 38433 10697 38669
rect 10933 38433 11023 38669
rect 11259 38433 11349 38669
rect 11585 38433 11675 38669
rect 11911 38433 12001 38669
rect 12237 38433 12327 38669
rect 12563 38433 12653 38669
rect 12889 38433 12979 38669
rect 13215 38433 13305 38669
rect 13541 38433 13631 38669
rect 13867 38433 13957 38669
rect 14193 38433 14283 38669
rect 14519 38433 14609 38669
rect 14845 38433 15000 38669
rect 0 38345 4967 38433
rect 9991 38345 15000 38433
rect 0 38109 241 38345
rect 477 38109 568 38345
rect 804 38109 895 38345
rect 1131 38109 1222 38345
rect 1458 38109 1549 38345
rect 1785 38109 1876 38345
rect 2112 38109 2203 38345
rect 2439 38109 2530 38345
rect 2766 38109 2857 38345
rect 3093 38109 3184 38345
rect 3420 38109 3511 38345
rect 3747 38109 3838 38345
rect 4074 38109 4165 38345
rect 4401 38109 4492 38345
rect 4728 38109 4819 38345
rect 9991 38109 10045 38345
rect 10281 38109 10371 38345
rect 10607 38109 10697 38345
rect 10933 38109 11023 38345
rect 11259 38109 11349 38345
rect 11585 38109 11675 38345
rect 11911 38109 12001 38345
rect 12237 38109 12327 38345
rect 12563 38109 12653 38345
rect 12889 38109 12979 38345
rect 13215 38109 13305 38345
rect 13541 38109 13631 38345
rect 13867 38109 13957 38345
rect 14193 38109 14283 38345
rect 14519 38109 14609 38345
rect 14845 38109 15000 38345
rect 0 38021 4967 38109
rect 9991 38021 15000 38109
rect 0 37785 241 38021
rect 477 37785 568 38021
rect 804 37785 895 38021
rect 1131 37785 1222 38021
rect 1458 37785 1549 38021
rect 1785 37785 1876 38021
rect 2112 37785 2203 38021
rect 2439 37785 2530 38021
rect 2766 37785 2857 38021
rect 3093 37785 3184 38021
rect 3420 37785 3511 38021
rect 3747 37785 3838 38021
rect 4074 37785 4165 38021
rect 4401 37785 4492 38021
rect 4728 37785 4819 38021
rect 9991 37785 10045 38021
rect 10281 37785 10371 38021
rect 10607 37785 10697 38021
rect 10933 37785 11023 38021
rect 11259 37785 11349 38021
rect 11585 37785 11675 38021
rect 11911 37785 12001 38021
rect 12237 37785 12327 38021
rect 12563 37785 12653 38021
rect 12889 37785 12979 38021
rect 13215 37785 13305 38021
rect 13541 37785 13631 38021
rect 13867 37785 13957 38021
rect 14193 37785 14283 38021
rect 14519 37785 14609 38021
rect 14845 37785 15000 38021
rect 0 37697 4967 37785
rect 9991 37697 15000 37785
rect 0 37461 241 37697
rect 477 37461 568 37697
rect 804 37461 895 37697
rect 1131 37461 1222 37697
rect 1458 37461 1549 37697
rect 1785 37461 1876 37697
rect 2112 37461 2203 37697
rect 2439 37461 2530 37697
rect 2766 37461 2857 37697
rect 3093 37461 3184 37697
rect 3420 37461 3511 37697
rect 3747 37461 3838 37697
rect 4074 37461 4165 37697
rect 4401 37461 4492 37697
rect 4728 37461 4819 37697
rect 9991 37461 10045 37697
rect 10281 37461 10371 37697
rect 10607 37461 10697 37697
rect 10933 37461 11023 37697
rect 11259 37461 11349 37697
rect 11585 37461 11675 37697
rect 11911 37461 12001 37697
rect 12237 37461 12327 37697
rect 12563 37461 12653 37697
rect 12889 37461 12979 37697
rect 13215 37461 13305 37697
rect 13541 37461 13631 37697
rect 13867 37461 13957 37697
rect 14193 37461 14283 37697
rect 14519 37461 14609 37697
rect 14845 37461 15000 37697
rect 0 37373 4967 37461
rect 9991 37373 15000 37461
rect 0 37137 241 37373
rect 477 37137 568 37373
rect 804 37137 895 37373
rect 1131 37198 1222 37373
rect 1458 37198 1549 37373
rect 1785 37198 1876 37373
rect 2112 37198 2203 37373
rect 2143 37137 2203 37198
rect 2439 37137 2530 37373
rect 2766 37137 2857 37373
rect 3093 37137 3184 37373
rect 3420 37137 3511 37373
rect 3747 37137 3838 37373
rect 4074 37137 4165 37373
rect 4401 37137 4492 37373
rect 4728 37137 4819 37373
rect 9991 37137 10045 37373
rect 10281 37137 10371 37373
rect 10607 37137 10697 37373
rect 10933 37137 11023 37373
rect 11259 37137 11349 37373
rect 11585 37137 11675 37373
rect 11911 37137 12001 37373
rect 12237 37137 12327 37373
rect 12563 37137 12653 37373
rect 12889 37195 12979 37373
rect 13215 37195 13305 37373
rect 13541 37195 13631 37373
rect 13867 37195 13957 37373
rect 14193 37137 14283 37373
rect 14519 37137 14609 37373
rect 14845 37137 15000 37373
rect 0 37049 959 37137
rect 2143 37049 4967 37137
rect 9991 37049 12823 37137
rect 14007 37049 15000 37137
rect 0 36813 241 37049
rect 477 36813 568 37049
rect 804 36813 895 37049
rect 2143 36813 2203 37049
rect 2439 36813 2530 37049
rect 2766 36813 2857 37049
rect 3093 36813 3184 37049
rect 3420 36813 3511 37049
rect 3747 36813 3838 37049
rect 4074 36813 4165 37049
rect 4401 36813 4492 37049
rect 4728 36813 4819 37049
rect 9991 36813 10045 37049
rect 10281 36813 10371 37049
rect 10607 36813 10697 37049
rect 10933 36813 11023 37049
rect 11259 36813 11349 37049
rect 11585 36813 11675 37049
rect 11911 36813 12001 37049
rect 12237 36813 12327 37049
rect 12563 36813 12653 37049
rect 14193 36813 14283 37049
rect 14519 36813 14609 37049
rect 14845 36813 15000 37049
rect 0 36725 959 36813
rect 2143 36725 4967 36813
rect 9991 36725 12823 36813
rect 14007 36725 15000 36813
rect 0 36489 241 36725
rect 477 36489 568 36725
rect 804 36489 895 36725
rect 2143 36494 2203 36725
rect 1131 36489 1222 36494
rect 1458 36489 1549 36494
rect 1785 36489 1876 36494
rect 2112 36489 2203 36494
rect 2439 36489 2530 36725
rect 2766 36489 2857 36725
rect 3093 36489 3184 36725
rect 3420 36489 3511 36725
rect 3747 36489 3838 36725
rect 4074 36489 4165 36725
rect 4401 36489 4492 36725
rect 4728 36489 4819 36725
rect 9991 36489 10045 36725
rect 10281 36489 10371 36725
rect 10607 36489 10697 36725
rect 10933 36489 11023 36725
rect 11259 36489 11349 36725
rect 11585 36489 11675 36725
rect 11911 36489 12001 36725
rect 12237 36489 12327 36725
rect 12563 36489 12653 36725
rect 12889 36489 12979 36491
rect 13215 36489 13305 36491
rect 13541 36489 13631 36491
rect 13867 36489 13957 36491
rect 14193 36489 14283 36725
rect 14519 36489 14609 36725
rect 14845 36489 15000 36725
rect 0 36401 4967 36489
rect 9991 36401 15000 36489
rect 0 36165 241 36401
rect 477 36165 568 36401
rect 804 36165 895 36401
rect 1131 36165 1222 36401
rect 1458 36165 1549 36401
rect 1785 36165 1876 36401
rect 2112 36165 2203 36401
rect 2439 36165 2530 36401
rect 2766 36165 2857 36401
rect 3093 36165 3184 36401
rect 3420 36165 3511 36401
rect 3747 36165 3838 36401
rect 4074 36165 4165 36401
rect 4401 36165 4492 36401
rect 4728 36165 4819 36401
rect 9991 36165 10045 36401
rect 10281 36165 10371 36401
rect 10607 36165 10697 36401
rect 10933 36165 11023 36401
rect 11259 36165 11349 36401
rect 11585 36165 11675 36401
rect 11911 36165 12001 36401
rect 12237 36165 12327 36401
rect 12563 36165 12653 36401
rect 12889 36165 12979 36401
rect 13215 36165 13305 36401
rect 13541 36165 13631 36401
rect 13867 36165 13957 36401
rect 14193 36165 14283 36401
rect 14519 36165 14609 36401
rect 14845 36165 15000 36401
rect 0 36077 4967 36165
rect 9991 36077 15000 36165
rect 0 35841 241 36077
rect 477 35841 568 36077
rect 804 35841 895 36077
rect 1131 35841 1222 36077
rect 1458 35841 1549 36077
rect 1785 35841 1876 36077
rect 2112 35841 2203 36077
rect 2439 35841 2530 36077
rect 2766 35841 2857 36077
rect 3093 35841 3184 36077
rect 3420 35841 3511 36077
rect 3747 35841 3838 36077
rect 4074 35841 4165 36077
rect 4401 35841 4492 36077
rect 4728 35841 4819 36077
rect 9991 35841 10045 36077
rect 10281 35841 10371 36077
rect 10607 35841 10697 36077
rect 10933 35841 11023 36077
rect 11259 35841 11349 36077
rect 11585 35841 11675 36077
rect 11911 35841 12001 36077
rect 12237 35841 12327 36077
rect 12563 35841 12653 36077
rect 12889 35841 12979 36077
rect 13215 35841 13305 36077
rect 13541 35841 13631 36077
rect 13867 35841 13957 36077
rect 14193 35841 14283 36077
rect 14519 35841 14609 36077
rect 14845 35841 15000 36077
rect 0 35753 4967 35841
rect 9991 35753 15000 35841
rect 0 35517 241 35753
rect 477 35517 568 35753
rect 804 35517 895 35753
rect 1131 35517 1222 35753
rect 1458 35517 1549 35753
rect 1785 35517 1876 35753
rect 2112 35517 2203 35753
rect 2439 35517 2530 35753
rect 2766 35517 2857 35753
rect 3093 35517 3184 35753
rect 3420 35517 3511 35753
rect 3747 35517 3838 35753
rect 4074 35517 4165 35753
rect 4401 35517 4492 35753
rect 4728 35517 4819 35753
rect 9991 35517 10045 35753
rect 10281 35517 10371 35753
rect 10607 35517 10697 35753
rect 10933 35517 11023 35753
rect 11259 35517 11349 35753
rect 11585 35517 11675 35753
rect 11911 35517 12001 35753
rect 12237 35517 12327 35753
rect 12563 35517 12653 35753
rect 12889 35517 12979 35753
rect 13215 35517 13305 35753
rect 13541 35517 13631 35753
rect 13867 35517 13957 35753
rect 14193 35517 14283 35753
rect 14519 35517 14609 35753
rect 14845 35517 15000 35753
rect 0 35429 4967 35517
rect 9991 35429 15000 35517
rect 0 35193 241 35429
rect 477 35193 568 35429
rect 804 35193 895 35429
rect 1131 35193 1222 35429
rect 1458 35193 1549 35429
rect 1785 35193 1876 35429
rect 2112 35193 2203 35429
rect 2439 35193 2530 35429
rect 2766 35193 2857 35429
rect 3093 35193 3184 35429
rect 3420 35193 3511 35429
rect 3747 35193 3838 35429
rect 4074 35193 4165 35429
rect 4401 35193 4492 35429
rect 4728 35193 4819 35429
rect 9991 35324 10045 35429
rect 5055 35193 5146 35324
rect 5382 35193 5473 35324
rect 5709 35193 5800 35324
rect 6036 35193 6127 35324
rect 6363 35193 6454 35324
rect 6690 35193 6781 35324
rect 7017 35193 7108 35324
rect 7344 35193 7435 35324
rect 7671 35193 7762 35324
rect 7998 35193 8089 35324
rect 8325 35193 8415 35324
rect 8651 35193 8741 35324
rect 8977 35193 9067 35324
rect 9303 35193 9393 35324
rect 9629 35193 9719 35324
rect 9955 35193 10045 35324
rect 10281 35193 10371 35429
rect 10607 35193 10697 35429
rect 10933 35193 11023 35429
rect 11259 35193 11349 35429
rect 11585 35193 11675 35429
rect 11911 35193 12001 35429
rect 12237 35193 12327 35429
rect 12563 35193 12653 35429
rect 12889 35193 12979 35429
rect 13215 35193 13305 35429
rect 13541 35193 13631 35429
rect 13867 35193 13957 35429
rect 14193 35193 14283 35429
rect 14519 35193 14609 35429
rect 14845 35193 15000 35429
rect 0 35157 15000 35193
tri 1933 34288 2265 34620 se
rect 2265 34596 12733 34620
tri 12733 34596 12757 34620 sw
rect 2265 34360 2268 34596
rect 2504 34588 2588 34596
rect 2824 34588 2908 34596
rect 3144 34360 3228 34596
rect 3464 34360 3548 34596
rect 3784 34360 3868 34596
rect 4104 34360 4188 34596
rect 4424 34360 4508 34596
rect 4744 34360 4828 34596
rect 5064 34360 5148 34596
rect 5384 34360 5468 34596
rect 5704 34360 5788 34596
rect 6024 34360 6108 34596
rect 6344 34360 6428 34596
rect 6664 34360 6748 34596
rect 6984 34360 7068 34596
rect 7304 34360 7388 34596
rect 7624 34360 7708 34596
rect 7944 34360 8028 34596
rect 8264 34360 8348 34596
rect 8584 34360 8668 34596
rect 8904 34360 8988 34596
rect 9224 34360 9308 34596
rect 9544 34360 9628 34596
rect 9864 34360 9948 34596
rect 10184 34360 10268 34596
rect 10504 34360 10588 34596
rect 10824 34360 10908 34596
rect 11144 34360 11228 34596
rect 11464 34360 11548 34596
rect 11784 34360 11868 34596
rect 12104 34587 12188 34596
rect 12424 34587 12508 34596
rect 12744 34360 12757 34596
rect 2265 34288 2331 34360
tri 1725 34080 1933 34288 se
rect 1933 34080 1946 34288
tri 1613 33968 1725 34080 se
rect 1725 34052 1946 34080
rect 2182 34124 2331 34288
rect 3035 34124 11961 34360
rect 2182 34123 11961 34124
rect 12665 34234 12757 34360
tri 12757 34234 13119 34596 sw
rect 12665 34123 12870 34234
rect 2182 34080 12870 34123
rect 2182 34052 2377 34080
rect 1725 33968 2377 34052
tri 2377 33968 2489 34080 nw
tri 1499 33854 1613 33968 se
rect 1613 33854 1626 33968
tri 1293 33648 1499 33854 se
rect 1499 33732 1626 33854
rect 1862 33732 2141 33968
tri 2141 33732 2377 33968 nw
tri 12509 33732 12857 34080 ne
rect 12857 33998 12870 34080
rect 13106 33998 13119 34234
rect 12857 33914 13119 33998
tri 13119 33914 13439 34234 sw
rect 12857 33732 13190 33914
rect 1499 33648 1725 33732
tri 970 33325 1293 33648 se
rect 1293 33412 1306 33648
rect 1542 33412 1725 33648
rect 1293 33325 1725 33412
tri 959 33314 970 33325 se
rect 970 33314 983 33325
rect 959 33089 983 33314
rect 1219 33316 1725 33325
tri 1725 33316 2141 33732 nw
tri 12857 33678 12911 33732 ne
rect 12911 33678 13190 33732
rect 13426 33678 13439 33914
tri 12911 33316 13273 33678 ne
rect 13273 33594 13439 33678
tri 13439 33594 13759 33914 sw
rect 13273 33358 13510 33594
rect 13746 33358 13759 33594
rect 13273 33316 13759 33358
rect 1219 33089 1499 33316
tri 1499 33090 1725 33316 nw
tri 13273 33090 13499 33316 ne
rect 13499 33314 13759 33316
tri 13759 33314 14039 33594 sw
rect 13499 33231 14039 33314
rect 959 33005 1499 33089
rect 959 32769 983 33005
rect 1219 32974 1499 33005
rect 959 32685 1035 32769
rect 959 32449 983 32685
rect 959 32365 1035 32449
rect 959 32129 983 32365
rect 959 32045 1035 32129
rect 959 31809 983 32045
rect 959 31725 1035 31809
rect 959 31489 983 31725
rect 959 31405 1035 31489
rect 959 31169 983 31405
rect 959 31085 1035 31169
rect 959 30849 983 31085
rect 959 30765 1035 30849
rect 959 30529 983 30765
rect 959 30445 1035 30529
rect 959 30209 983 30445
rect 959 30125 1035 30209
rect 959 29889 983 30125
rect 959 29805 1035 29889
rect 959 29569 983 29805
rect 959 29485 1035 29569
rect 959 29249 983 29485
rect 959 29165 1035 29249
rect 959 28929 983 29165
rect 959 28845 1035 28929
rect 959 28609 983 28845
rect 959 28525 1035 28609
rect 959 28289 983 28525
rect 959 28205 1035 28289
rect 959 27969 983 28205
rect 959 27885 1035 27969
rect 959 27649 983 27885
rect 959 27565 1035 27649
rect 959 27329 983 27565
rect 959 27245 1035 27329
rect 959 27009 983 27245
rect 959 26925 1035 27009
rect 959 26689 983 26925
rect 959 26605 1035 26689
rect 959 26369 983 26605
rect 959 26285 1035 26369
rect 959 26049 983 26285
rect 959 25965 1035 26049
rect 959 25729 983 25965
rect 959 25645 1035 25729
rect 959 25409 983 25645
rect 959 25325 1035 25409
rect 959 25089 983 25325
rect 959 25005 1035 25089
rect 959 24769 983 25005
rect 959 24685 1035 24769
rect 959 24449 983 24685
rect 959 24365 1035 24449
rect 959 24129 983 24365
rect 959 24045 1035 24129
rect 959 23809 983 24045
rect 959 23725 1035 23809
rect 959 23489 983 23725
rect 959 23405 1035 23489
rect 959 23169 983 23405
rect 959 23085 1035 23169
rect 959 22849 983 23085
rect 959 22765 1035 22849
rect 959 22529 983 22765
rect 959 22445 1035 22529
rect 959 22209 983 22445
rect 959 22125 1035 22209
rect 959 21889 983 22125
rect 959 21805 1035 21889
rect 959 21569 983 21805
rect 959 21485 1035 21569
rect 959 21249 983 21485
rect 959 21230 1035 21249
rect 1419 21230 1499 32974
rect 959 21165 1499 21230
rect 959 20929 983 21165
rect 1219 20929 1499 21165
rect 13499 32995 13779 33231
rect 14015 32995 14039 33231
rect 13499 32911 14039 32995
rect 13499 32866 13779 32911
rect 13499 21122 13581 32866
rect 14015 32675 14039 32911
rect 13965 32591 14039 32675
rect 14015 32355 14039 32591
rect 13965 32271 14039 32355
rect 14015 32035 14039 32271
rect 13965 31951 14039 32035
rect 14015 31715 14039 31951
rect 13965 31631 14039 31715
rect 14015 31395 14039 31631
rect 13965 31311 14039 31395
rect 14015 31075 14039 31311
rect 13965 30991 14039 31075
rect 14015 30755 14039 30991
rect 13965 30671 14039 30755
rect 14015 30435 14039 30671
rect 13965 30351 14039 30435
rect 14015 30115 14039 30351
rect 13965 30031 14039 30115
rect 14015 29795 14039 30031
rect 13965 29711 14039 29795
rect 14015 29475 14039 29711
rect 13965 29391 14039 29475
rect 14015 29155 14039 29391
rect 13965 29071 14039 29155
rect 14015 28835 14039 29071
rect 13965 28751 14039 28835
rect 14015 28515 14039 28751
rect 13965 28431 14039 28515
rect 14015 28195 14039 28431
rect 13965 28111 14039 28195
rect 14015 27875 14039 28111
rect 13965 27791 14039 27875
rect 14015 27555 14039 27791
rect 13965 27471 14039 27555
rect 14015 27235 14039 27471
rect 13965 27151 14039 27235
rect 14015 26915 14039 27151
rect 13965 26831 14039 26915
rect 14015 26595 14039 26831
rect 13965 26511 14039 26595
rect 14015 26275 14039 26511
rect 13965 26191 14039 26275
rect 14015 25955 14039 26191
rect 13965 25871 14039 25955
rect 14015 25635 14039 25871
rect 13965 25551 14039 25635
rect 14015 25315 14039 25551
rect 13965 25231 14039 25315
rect 14015 24995 14039 25231
rect 13965 24911 14039 24995
rect 14015 24675 14039 24911
rect 13965 24591 14039 24675
rect 14015 24355 14039 24591
rect 13965 24271 14039 24355
rect 14015 24035 14039 24271
rect 13965 23951 14039 24035
rect 14015 23715 14039 23951
rect 13965 23631 14039 23715
rect 14015 23395 14039 23631
rect 13965 23311 14039 23395
rect 14015 23075 14039 23311
rect 13965 22991 14039 23075
rect 14015 22755 14039 22991
rect 13965 22671 14039 22755
rect 14015 22435 14039 22671
rect 13965 22351 14039 22435
rect 14015 22115 14039 22351
rect 13965 22031 14039 22115
rect 14015 21795 14039 22031
rect 13965 21711 14039 21795
rect 14015 21475 14039 21711
rect 13965 21391 14039 21475
rect 14015 21155 14039 21391
rect 13965 21122 14039 21155
rect 13499 21071 14039 21122
rect 959 20846 1499 20929
tri 959 20566 1239 20846 ne
rect 1239 20802 1499 20846
rect 1239 20566 1252 20802
rect 1488 20566 1499 20802
tri 1239 20306 1499 20566 ne
tri 1499 20482 2087 21070 sw
tri 13273 20844 13499 21070 se
rect 13499 20844 13779 21071
rect 1499 20306 1572 20482
tri 1499 20246 1559 20306 ne
rect 1559 20246 1572 20306
rect 1808 20306 2087 20482
tri 2087 20306 2263 20482 sw
tri 12857 20428 13273 20844 se
rect 13273 20835 13779 20844
rect 14015 20846 14039 21071
rect 14015 20835 14028 20846
tri 14028 20835 14039 20846 nw
rect 13273 20748 13705 20835
rect 13273 20512 13456 20748
rect 13692 20512 13705 20748
tri 13705 20512 14028 20835 nw
rect 13273 20428 13385 20512
tri 12735 20306 12857 20428 se
rect 12857 20306 13136 20428
rect 1808 20246 2263 20306
tri 1559 19926 1879 20246 ne
rect 1879 20162 2263 20246
rect 1879 19926 1892 20162
rect 2128 20080 2263 20162
tri 2263 20080 2489 20306 sw
tri 12509 20080 12735 20306 se
rect 12735 20192 13136 20306
rect 13372 20192 13385 20428
tri 13385 20192 13705 20512 nw
rect 12735 20108 13065 20192
rect 12735 20080 12816 20108
rect 2128 20040 12816 20080
rect 2128 19926 2308 20040
tri 1879 19564 2241 19926 ne
rect 2241 19800 2308 19926
rect 12692 19872 12816 20040
rect 13052 19872 13065 20108
tri 13065 19872 13385 20192 nw
rect 12692 19800 12733 19872
rect 2241 19564 2254 19800
rect 2490 19564 2574 19576
rect 2810 19564 2894 19576
rect 3130 19564 3214 19576
rect 3450 19564 3534 19576
rect 3770 19564 3854 19576
rect 4090 19564 4174 19576
rect 4410 19564 4494 19576
rect 4730 19564 4814 19576
rect 5050 19564 5134 19576
rect 5370 19564 5454 19576
rect 5690 19564 5774 19576
rect 6010 19564 6094 19576
rect 6330 19564 6414 19576
rect 6650 19564 6734 19576
rect 6970 19564 7054 19576
rect 7290 19564 7374 19576
rect 7610 19564 7694 19576
rect 7930 19564 8014 19576
rect 8250 19564 8334 19576
rect 8570 19564 8654 19576
rect 8890 19564 8974 19576
rect 9210 19564 9294 19576
rect 9530 19564 9614 19576
rect 9850 19564 9934 19576
rect 10170 19564 10254 19576
rect 10490 19564 10574 19576
rect 10810 19564 10894 19576
rect 11130 19564 11214 19576
rect 11450 19564 11534 19576
rect 11770 19564 11854 19576
rect 12090 19564 12174 19576
rect 12410 19564 12494 19576
rect 12730 19564 12733 19800
tri 2241 19540 2265 19564 ne
rect 2265 19540 12733 19564
tri 12733 19540 13065 19872 nw
tri 6504 19140 6904 19540 ne
rect 0 18972 5622 19000
rect 0 18736 143 18972
rect 379 18736 465 18972
rect 701 18736 787 18972
rect 1023 18736 1109 18972
rect 1345 18736 1431 18972
rect 1667 18736 1753 18972
rect 1989 18736 2075 18972
rect 2311 18736 2397 18972
rect 2633 18736 2719 18972
rect 2955 18908 3041 18972
rect 3277 18908 3363 18972
rect 3599 18908 3685 18972
rect 3921 18908 4007 18972
rect 4243 18908 4329 18972
rect 4565 18908 4651 18972
rect 4887 18908 4973 18972
rect 5209 18908 5295 18972
rect 5234 18736 5295 18908
rect 5531 18800 5622 18972
tri 5622 18800 5822 19000 sw
rect 5531 18736 5822 18800
rect 0 18636 2930 18736
rect 5234 18636 5822 18736
rect 0 18400 143 18636
rect 379 18400 465 18636
rect 701 18400 787 18636
rect 1023 18400 1109 18636
rect 1345 18400 1431 18636
rect 1667 18400 1753 18636
rect 1989 18400 2075 18636
rect 2311 18400 2397 18636
rect 2633 18400 2719 18636
rect 5234 18400 5295 18636
rect 5531 18400 5822 18636
rect 0 18300 2930 18400
rect 5234 18300 5822 18400
rect 0 18064 143 18300
rect 379 18064 465 18300
rect 701 18064 787 18300
rect 1023 18064 1109 18300
rect 1345 18064 1431 18300
rect 1667 18064 1753 18300
rect 1989 18064 2075 18300
rect 2311 18064 2397 18300
rect 2633 18064 2719 18300
rect 5234 18064 5295 18300
rect 5531 18064 5822 18300
rect 0 17964 2930 18064
rect 5234 17964 5822 18064
rect 0 17728 143 17964
rect 379 17728 465 17964
rect 701 17728 787 17964
rect 1023 17728 1109 17964
rect 1345 17728 1431 17964
rect 1667 17728 1753 17964
rect 1989 17728 2075 17964
rect 2311 17728 2397 17964
rect 2633 17728 2719 17964
rect 5234 17728 5295 17964
rect 5531 17728 5822 17964
rect 0 17628 2930 17728
rect 5234 17628 5822 17728
rect 0 17392 143 17628
rect 379 17392 465 17628
rect 701 17392 787 17628
rect 1023 17392 1109 17628
rect 1345 17392 1431 17628
rect 1667 17392 1753 17628
rect 1989 17392 2075 17628
rect 2311 17392 2397 17628
rect 2633 17392 2719 17628
rect 5234 17392 5295 17628
rect 5531 17392 5822 17628
rect 0 17324 2930 17392
rect 5234 17324 5822 17392
rect 0 17292 5822 17324
rect 0 17056 143 17292
rect 379 17056 465 17292
rect 701 17056 787 17292
rect 1023 17056 1109 17292
rect 1345 17056 1431 17292
rect 1667 17056 1753 17292
rect 1989 17056 2075 17292
rect 2311 17056 2397 17292
rect 2633 17056 2719 17292
rect 2955 17056 3041 17292
rect 3277 17231 3363 17292
rect 3599 17231 3685 17292
rect 3921 17231 4007 17292
rect 4243 17231 4329 17292
rect 4565 17231 4651 17292
rect 4887 17231 4973 17292
rect 5209 17231 5295 17292
rect 5235 17087 5295 17231
rect 3277 17056 3363 17087
rect 3599 17056 3685 17087
rect 3921 17056 4007 17087
rect 4243 17056 4329 17087
rect 4565 17056 4651 17087
rect 4887 17056 4973 17087
rect 5209 17056 5295 17087
rect 5531 17056 5822 17292
rect 0 16956 5822 17056
rect 0 16720 143 16956
rect 379 16720 465 16956
rect 701 16720 787 16956
rect 1023 16720 1109 16956
rect 1345 16720 1431 16956
rect 1667 16720 1753 16956
rect 1989 16720 2075 16956
rect 2311 16720 2397 16956
rect 2633 16720 2719 16956
rect 2955 16720 3041 16956
rect 3277 16720 3363 16956
rect 3599 16720 3685 16956
rect 3921 16720 4007 16956
rect 4243 16720 4329 16956
rect 4565 16720 4651 16956
rect 4887 16720 4973 16956
rect 5209 16720 5295 16956
rect 5531 16720 5822 16956
rect 0 16620 5822 16720
rect 0 16384 143 16620
rect 379 16384 465 16620
rect 701 16384 787 16620
rect 1023 16384 1109 16620
rect 1345 16384 1431 16620
rect 1667 16384 1753 16620
rect 1989 16384 2075 16620
rect 2311 16384 2397 16620
rect 2633 16384 2719 16620
rect 2955 16384 3041 16620
rect 3277 16384 3363 16620
rect 3599 16384 3685 16620
rect 3921 16384 4007 16620
rect 4243 16384 4329 16620
rect 4565 16384 4651 16620
rect 4887 16384 4973 16620
rect 5209 16384 5295 16620
rect 5531 16384 5822 16620
rect 0 16284 5822 16384
rect 0 16048 143 16284
rect 379 16048 465 16284
rect 701 16048 787 16284
rect 1023 16048 1109 16284
rect 1345 16048 1431 16284
rect 1667 16048 1753 16284
rect 1989 16048 2075 16284
rect 2311 16048 2397 16284
rect 2633 16048 2719 16284
rect 2955 16048 3041 16284
rect 3277 16048 3363 16284
rect 3599 16048 3685 16284
rect 3921 16048 4007 16284
rect 4243 16048 4329 16284
rect 4565 16048 4651 16284
rect 4887 16048 4973 16284
rect 5209 16048 5295 16284
rect 5531 16048 5822 16284
rect 0 15948 5822 16048
rect 0 15712 143 15948
rect 379 15712 465 15948
rect 701 15712 787 15948
rect 1023 15712 1109 15948
rect 1345 15712 1431 15948
rect 1667 15712 1753 15948
rect 1989 15712 2075 15948
rect 2311 15712 2397 15948
rect 2633 15712 2719 15948
rect 2955 15712 3041 15948
rect 3277 15712 3363 15948
rect 3599 15712 3685 15948
rect 3921 15712 4007 15948
rect 4243 15712 4329 15948
rect 4565 15712 4651 15948
rect 4887 15712 4973 15948
rect 5209 15712 5295 15948
rect 5531 15712 5822 15948
rect 0 15612 5822 15712
rect 0 15376 143 15612
rect 379 15376 465 15612
rect 701 15376 787 15612
rect 1023 15376 1109 15612
rect 1345 15376 1431 15612
rect 1667 15376 1753 15612
rect 1989 15376 2075 15612
rect 2311 15376 2397 15612
rect 2633 15376 2719 15612
rect 2955 15376 3041 15612
rect 3277 15376 3363 15612
rect 3599 15376 3685 15612
rect 3921 15376 4007 15612
rect 4243 15376 4329 15612
rect 4565 15376 4651 15612
rect 4887 15376 4973 15612
rect 5209 15376 5295 15612
rect 5531 15376 5822 15612
rect 0 15276 5822 15376
rect 0 15040 143 15276
rect 379 15040 465 15276
rect 701 15040 787 15276
rect 1023 15040 1109 15276
rect 1345 15040 1431 15276
rect 1667 15040 1753 15276
rect 1989 15040 2075 15276
rect 2311 15040 2397 15276
rect 2633 15040 2719 15276
rect 2955 15040 3041 15276
rect 3277 15040 3363 15276
rect 3599 15040 3685 15276
rect 3921 15040 4007 15276
rect 4243 15040 4329 15276
rect 4565 15040 4651 15276
rect 4887 15040 4973 15276
rect 5209 15040 5295 15276
rect 5531 15040 5822 15276
rect 0 14940 5822 15040
rect 0 14704 143 14940
rect 379 14704 465 14940
rect 701 14704 787 14940
rect 1023 14718 1109 14940
rect 1345 14718 1431 14940
rect 1667 14718 1753 14940
rect 1989 14718 2075 14940
rect 2022 14704 2075 14718
rect 2311 14704 2397 14940
rect 2633 14704 2719 14940
rect 2955 14704 3041 14940
rect 3277 14704 3363 14940
rect 3599 14704 3685 14940
rect 3921 14704 4007 14940
rect 4243 14704 4329 14940
rect 4565 14704 4651 14940
rect 4887 14704 4973 14940
rect 5209 14704 5295 14940
rect 5531 14704 5822 14940
rect 0 14604 918 14704
rect 2022 14604 5822 14704
rect 0 14368 143 14604
rect 379 14368 465 14604
rect 701 14368 787 14604
rect 2022 14368 2075 14604
rect 2311 14368 2397 14604
rect 2633 14368 2719 14604
rect 2955 14368 3041 14604
rect 3277 14368 3363 14604
rect 3599 14368 3685 14604
rect 3921 14368 4007 14604
rect 4243 14368 4329 14604
rect 4565 14368 4651 14604
rect 4887 14368 4973 14604
rect 5209 14368 5295 14604
rect 5531 14368 5822 14604
rect 0 14334 918 14368
rect 2022 14334 5822 14368
rect 0 14268 5822 14334
rect 0 14032 143 14268
rect 379 14032 465 14268
rect 701 14032 787 14268
rect 1023 14032 1109 14268
rect 1345 14032 1431 14268
rect 1667 14032 1753 14268
rect 1989 14032 2075 14268
rect 2311 14032 2397 14268
rect 2633 14032 2719 14268
rect 2955 14032 3041 14268
rect 3277 14032 3363 14268
rect 3599 14032 3685 14268
rect 3921 14032 4007 14268
rect 4243 14032 4329 14268
rect 4565 14032 4651 14268
rect 4887 14032 4973 14268
rect 5209 14032 5295 14268
rect 5531 14207 5822 14268
rect 5531 14032 5622 14207
rect 0 14007 5622 14032
tri 5622 14007 5822 14207 nw
rect 6904 14009 8104 19540
tri 8104 19140 8504 19540 nw
tri 9140 18800 9340 19000 se
rect 9340 18972 15000 19000
rect 9340 18800 9469 18972
rect 9140 18736 9469 18800
rect 9705 18908 9790 18972
rect 10026 18908 10111 18972
rect 10347 18908 10432 18972
rect 10668 18908 10753 18972
rect 10989 18908 11074 18972
rect 11310 18908 11395 18972
rect 11631 18908 11716 18972
rect 11952 18908 12037 18972
rect 9705 18736 9730 18908
rect 12034 18736 12037 18908
rect 12273 18736 12358 18972
rect 12594 18736 12679 18972
rect 12915 18736 13000 18972
rect 13236 18736 13321 18972
rect 13557 18736 13642 18972
rect 13878 18736 13963 18972
rect 14199 18736 14284 18972
rect 14520 18736 14605 18972
rect 14841 18736 15000 18972
rect 9140 18636 9730 18736
rect 12034 18636 15000 18736
rect 9140 18400 9469 18636
rect 9705 18400 9730 18636
rect 12034 18400 12037 18636
rect 12273 18400 12358 18636
rect 12594 18400 12679 18636
rect 12915 18400 13000 18636
rect 13236 18400 13321 18636
rect 13557 18400 13642 18636
rect 13878 18400 13963 18636
rect 14199 18400 14284 18636
rect 14520 18400 14605 18636
rect 14841 18400 15000 18636
rect 9140 18300 9730 18400
rect 12034 18300 15000 18400
rect 9140 18064 9469 18300
rect 9705 18064 9730 18300
rect 12034 18064 12037 18300
rect 12273 18064 12358 18300
rect 12594 18064 12679 18300
rect 12915 18064 13000 18300
rect 13236 18064 13321 18300
rect 13557 18064 13642 18300
rect 13878 18064 13963 18300
rect 14199 18064 14284 18300
rect 14520 18064 14605 18300
rect 14841 18064 15000 18300
rect 9140 17964 9730 18064
rect 12034 17964 15000 18064
rect 9140 17728 9469 17964
rect 9705 17728 9730 17964
rect 12034 17728 12037 17964
rect 12273 17728 12358 17964
rect 12594 17728 12679 17964
rect 12915 17728 13000 17964
rect 13236 17728 13321 17964
rect 13557 17728 13642 17964
rect 13878 17728 13963 17964
rect 14199 17728 14284 17964
rect 14520 17728 14605 17964
rect 14841 17728 15000 17964
rect 9140 17628 9730 17728
rect 12034 17628 15000 17728
rect 9140 17392 9469 17628
rect 9705 17392 9730 17628
rect 12034 17392 12037 17628
rect 12273 17392 12358 17628
rect 12594 17392 12679 17628
rect 12915 17392 13000 17628
rect 13236 17392 13321 17628
rect 13557 17392 13642 17628
rect 13878 17392 13963 17628
rect 14199 17392 14284 17628
rect 14520 17392 14605 17628
rect 14841 17392 15000 17628
rect 9140 17324 9730 17392
rect 12034 17324 15000 17392
rect 9140 17292 15000 17324
rect 9140 17056 9469 17292
rect 9705 17231 9790 17292
rect 10026 17231 10111 17292
rect 10347 17231 10432 17292
rect 10668 17231 10753 17292
rect 10989 17231 11074 17292
rect 11310 17231 11395 17292
rect 11631 17231 11716 17292
rect 9705 17087 9727 17231
rect 9705 17056 9790 17087
rect 10026 17056 10111 17087
rect 10347 17056 10432 17087
rect 10668 17056 10753 17087
rect 10989 17056 11074 17087
rect 11310 17056 11395 17087
rect 11631 17056 11716 17087
rect 11952 17056 12037 17292
rect 12273 17056 12358 17292
rect 12594 17056 12679 17292
rect 12915 17056 13000 17292
rect 13236 17056 13321 17292
rect 13557 17056 13642 17292
rect 13878 17056 13963 17292
rect 14199 17056 14284 17292
rect 14520 17056 14605 17292
rect 14841 17056 15000 17292
rect 9140 16956 15000 17056
rect 9140 16720 9469 16956
rect 9705 16720 9790 16956
rect 10026 16720 10111 16956
rect 10347 16720 10432 16956
rect 10668 16720 10753 16956
rect 10989 16720 11074 16956
rect 11310 16720 11395 16956
rect 11631 16720 11716 16956
rect 11952 16720 12037 16956
rect 12273 16720 12358 16956
rect 12594 16720 12679 16956
rect 12915 16720 13000 16956
rect 13236 16720 13321 16956
rect 13557 16720 13642 16956
rect 13878 16720 13963 16956
rect 14199 16720 14284 16956
rect 14520 16720 14605 16956
rect 14841 16720 15000 16956
rect 9140 16620 15000 16720
rect 9140 16384 9469 16620
rect 9705 16384 9790 16620
rect 10026 16384 10111 16620
rect 10347 16384 10432 16620
rect 10668 16384 10753 16620
rect 10989 16384 11074 16620
rect 11310 16384 11395 16620
rect 11631 16384 11716 16620
rect 11952 16384 12037 16620
rect 12273 16384 12358 16620
rect 12594 16384 12679 16620
rect 12915 16384 13000 16620
rect 13236 16384 13321 16620
rect 13557 16384 13642 16620
rect 13878 16384 13963 16620
rect 14199 16384 14284 16620
rect 14520 16384 14605 16620
rect 14841 16384 15000 16620
rect 9140 16284 15000 16384
rect 9140 16048 9469 16284
rect 9705 16048 9790 16284
rect 10026 16048 10111 16284
rect 10347 16048 10432 16284
rect 10668 16048 10753 16284
rect 10989 16048 11074 16284
rect 11310 16048 11395 16284
rect 11631 16048 11716 16284
rect 11952 16048 12037 16284
rect 12273 16048 12358 16284
rect 12594 16048 12679 16284
rect 12915 16048 13000 16284
rect 13236 16048 13321 16284
rect 13557 16048 13642 16284
rect 13878 16048 13963 16284
rect 14199 16048 14284 16284
rect 14520 16048 14605 16284
rect 14841 16048 15000 16284
rect 9140 15948 15000 16048
rect 9140 15712 9469 15948
rect 9705 15712 9790 15948
rect 10026 15712 10111 15948
rect 10347 15712 10432 15948
rect 10668 15712 10753 15948
rect 10989 15712 11074 15948
rect 11310 15712 11395 15948
rect 11631 15712 11716 15948
rect 11952 15712 12037 15948
rect 12273 15712 12358 15948
rect 12594 15712 12679 15948
rect 12915 15712 13000 15948
rect 13236 15712 13321 15948
rect 13557 15712 13642 15948
rect 13878 15712 13963 15948
rect 14199 15712 14284 15948
rect 14520 15712 14605 15948
rect 14841 15712 15000 15948
rect 9140 15612 15000 15712
rect 9140 15376 9469 15612
rect 9705 15376 9790 15612
rect 10026 15376 10111 15612
rect 10347 15376 10432 15612
rect 10668 15376 10753 15612
rect 10989 15376 11074 15612
rect 11310 15376 11395 15612
rect 11631 15376 11716 15612
rect 11952 15376 12037 15612
rect 12273 15376 12358 15612
rect 12594 15376 12679 15612
rect 12915 15376 13000 15612
rect 13236 15376 13321 15612
rect 13557 15376 13642 15612
rect 13878 15376 13963 15612
rect 14199 15376 14284 15612
rect 14520 15376 14605 15612
rect 14841 15376 15000 15612
rect 9140 15276 15000 15376
rect 9140 15040 9469 15276
rect 9705 15040 9790 15276
rect 10026 15040 10111 15276
rect 10347 15040 10432 15276
rect 10668 15040 10753 15276
rect 10989 15040 11074 15276
rect 11310 15040 11395 15276
rect 11631 15040 11716 15276
rect 11952 15040 12037 15276
rect 12273 15040 12358 15276
rect 12594 15040 12679 15276
rect 12915 15040 13000 15276
rect 13236 15040 13321 15276
rect 13557 15040 13642 15276
rect 13878 15040 13963 15276
rect 14199 15040 14284 15276
rect 14520 15040 14605 15276
rect 14841 15040 15000 15276
rect 9140 14940 15000 15040
rect 9140 14704 9469 14940
rect 9705 14704 9790 14940
rect 10026 14704 10111 14940
rect 10347 14704 10432 14940
rect 10668 14704 10753 14940
rect 10989 14704 11074 14940
rect 11310 14704 11395 14940
rect 11631 14704 11716 14940
rect 11952 14704 12037 14940
rect 12273 14704 12358 14940
rect 12594 14704 12679 14940
rect 12915 14718 13000 14940
rect 13236 14718 13321 14940
rect 13557 14718 13642 14940
rect 13878 14718 13963 14940
rect 12915 14704 12918 14718
rect 14199 14704 14284 14940
rect 14520 14704 14605 14940
rect 14841 14704 15000 14940
rect 9140 14604 12918 14704
rect 14022 14604 15000 14704
rect 9140 14368 9469 14604
rect 9705 14368 9790 14604
rect 10026 14368 10111 14604
rect 10347 14368 10432 14604
rect 10668 14368 10753 14604
rect 10989 14368 11074 14604
rect 11310 14368 11395 14604
rect 11631 14368 11716 14604
rect 11952 14368 12037 14604
rect 12273 14368 12358 14604
rect 12594 14368 12679 14604
rect 12915 14368 12918 14604
rect 14199 14368 14284 14604
rect 14520 14368 14605 14604
rect 14841 14368 15000 14604
rect 9140 14334 12918 14368
rect 14022 14334 15000 14368
rect 9140 14268 15000 14334
rect 9140 14207 9469 14268
tri 9140 14007 9340 14207 ne
rect 9340 14032 9469 14207
rect 9705 14032 9790 14268
rect 10026 14032 10111 14268
rect 10347 14032 10432 14268
rect 10668 14032 10753 14268
rect 10989 14032 11074 14268
rect 11310 14032 11395 14268
rect 11631 14032 11716 14268
rect 11952 14032 12037 14268
rect 12273 14032 12358 14268
rect 12594 14032 12679 14268
rect 12915 14032 13000 14268
rect 13236 14032 13321 14268
rect 13557 14032 13642 14268
rect 13878 14032 13963 14268
rect 14199 14032 14284 14268
rect 14520 14032 14605 14268
rect 14841 14032 15000 14268
rect 9340 14007 15000 14032
<< via4 >>
rect 241 39729 477 39965
rect 568 39729 804 39965
rect 895 39729 1131 39965
rect 1222 39729 1458 39965
rect 1549 39729 1785 39965
rect 1876 39729 2112 39965
rect 2203 39729 2439 39965
rect 2530 39729 2766 39965
rect 2857 39729 3093 39965
rect 3184 39729 3420 39965
rect 3511 39729 3747 39965
rect 3838 39729 4074 39965
rect 4165 39729 4401 39965
rect 4492 39729 4728 39965
rect 4819 39729 5055 39965
rect 5146 39870 5382 39965
rect 5473 39870 5709 39965
rect 5800 39870 6036 39965
rect 6127 39870 6363 39965
rect 6454 39870 6690 39965
rect 6781 39870 7017 39965
rect 7108 39870 7344 39965
rect 7435 39870 7671 39965
rect 7762 39870 7998 39965
rect 8089 39870 8325 39965
rect 8415 39870 8651 39965
rect 8741 39870 8977 39965
rect 9067 39870 9303 39965
rect 9393 39870 9629 39965
rect 9719 39870 9955 39965
rect 5146 39729 5259 39870
rect 5259 39729 5382 39870
rect 5473 39729 5709 39870
rect 5800 39729 6036 39870
rect 6127 39729 6363 39870
rect 6454 39729 6690 39870
rect 6781 39729 7017 39870
rect 7108 39729 7344 39870
rect 7435 39729 7671 39870
rect 7762 39729 7998 39870
rect 8089 39729 8325 39870
rect 8415 39729 8651 39870
rect 8741 39729 8977 39870
rect 9067 39729 9303 39870
rect 9393 39729 9629 39870
rect 9719 39729 9723 39870
rect 9723 39729 9955 39870
rect 10045 39729 10281 39965
rect 10371 39729 10607 39965
rect 10697 39729 10933 39965
rect 11023 39729 11259 39965
rect 11349 39729 11585 39965
rect 11675 39729 11911 39965
rect 12001 39729 12237 39965
rect 12327 39729 12563 39965
rect 12653 39729 12889 39965
rect 12979 39729 13215 39965
rect 13305 39729 13541 39965
rect 13631 39729 13867 39965
rect 13957 39729 14193 39965
rect 14283 39729 14519 39965
rect 14609 39729 14845 39965
rect 241 39405 477 39641
rect 568 39405 804 39641
rect 895 39405 1131 39641
rect 1222 39405 1458 39641
rect 1549 39405 1785 39641
rect 1876 39405 2112 39641
rect 2203 39405 2439 39641
rect 2530 39405 2766 39641
rect 2857 39405 3093 39641
rect 3184 39405 3420 39641
rect 3511 39405 3747 39641
rect 3838 39405 4074 39641
rect 4165 39405 4401 39641
rect 4492 39405 4728 39641
rect 4819 39468 5055 39641
rect 5146 39566 5259 39641
rect 5259 39566 5382 39641
rect 5473 39566 5709 39641
rect 5800 39566 6036 39641
rect 6127 39566 6363 39641
rect 6454 39566 6690 39641
rect 6781 39566 7017 39641
rect 7108 39566 7344 39641
rect 7435 39566 7671 39641
rect 7762 39566 7998 39641
rect 8089 39566 8325 39641
rect 8415 39566 8651 39641
rect 8741 39566 8977 39641
rect 9067 39566 9303 39641
rect 9393 39566 9629 39641
rect 9719 39566 9723 39641
rect 9723 39566 9955 39641
rect 5146 39468 5382 39566
rect 5473 39468 5709 39566
rect 5800 39468 6036 39566
rect 6127 39468 6363 39566
rect 6454 39468 6690 39566
rect 6781 39468 7017 39566
rect 7108 39468 7344 39566
rect 7435 39468 7671 39566
rect 7762 39468 7998 39566
rect 8089 39468 8325 39566
rect 8415 39468 8651 39566
rect 8741 39468 8977 39566
rect 9067 39468 9303 39566
rect 9393 39468 9629 39566
rect 9719 39468 9955 39566
rect 4819 39405 4967 39468
rect 4967 39405 5055 39468
rect 5146 39405 5382 39468
rect 5473 39405 5709 39468
rect 5800 39405 6036 39468
rect 6127 39405 6363 39468
rect 6454 39405 6690 39468
rect 6781 39405 7017 39468
rect 7108 39405 7344 39468
rect 7435 39405 7671 39468
rect 7762 39405 7998 39468
rect 8089 39405 8325 39468
rect 8415 39405 8651 39468
rect 8741 39405 8977 39468
rect 9067 39405 9303 39468
rect 9393 39405 9629 39468
rect 9719 39405 9955 39468
rect 10045 39405 10281 39641
rect 10371 39405 10607 39641
rect 10697 39405 10933 39641
rect 11023 39405 11259 39641
rect 11349 39405 11585 39641
rect 11675 39405 11911 39641
rect 12001 39405 12237 39641
rect 12327 39405 12563 39641
rect 12653 39405 12889 39641
rect 12979 39405 13215 39641
rect 13305 39405 13541 39641
rect 13631 39405 13867 39641
rect 13957 39405 14193 39641
rect 14283 39405 14519 39641
rect 14609 39405 14845 39641
rect 241 39081 477 39317
rect 568 39081 804 39317
rect 895 39081 1131 39317
rect 1222 39081 1458 39317
rect 1549 39081 1785 39317
rect 1876 39081 2112 39317
rect 2203 39081 2439 39317
rect 2530 39081 2766 39317
rect 2857 39081 3093 39317
rect 3184 39081 3420 39317
rect 3511 39081 3747 39317
rect 3838 39081 4074 39317
rect 4165 39081 4401 39317
rect 4492 39081 4728 39317
rect 4819 39081 4967 39317
rect 4967 39081 5055 39317
rect 5146 39081 5382 39317
rect 5473 39081 5709 39317
rect 5800 39081 6036 39317
rect 6127 39081 6363 39317
rect 6454 39081 6690 39317
rect 6781 39081 7017 39317
rect 7108 39081 7344 39317
rect 7435 39081 7671 39317
rect 7762 39081 7998 39317
rect 8089 39081 8325 39317
rect 8415 39081 8651 39317
rect 8741 39081 8977 39317
rect 9067 39081 9303 39317
rect 9393 39081 9629 39317
rect 9719 39081 9955 39317
rect 10045 39081 10281 39317
rect 10371 39081 10607 39317
rect 10697 39081 10933 39317
rect 11023 39081 11259 39317
rect 11349 39081 11585 39317
rect 11675 39081 11911 39317
rect 12001 39081 12237 39317
rect 12327 39081 12563 39317
rect 12653 39081 12889 39317
rect 12979 39081 13215 39317
rect 13305 39081 13541 39317
rect 13631 39081 13867 39317
rect 13957 39081 14193 39317
rect 14283 39081 14519 39317
rect 14609 39081 14845 39317
rect 241 38757 477 38993
rect 568 38757 804 38993
rect 895 38757 1131 38993
rect 1222 38757 1458 38993
rect 1549 38757 1785 38993
rect 1876 38757 2112 38993
rect 2203 38757 2439 38993
rect 2530 38757 2766 38993
rect 2857 38757 3093 38993
rect 3184 38757 3420 38993
rect 3511 38757 3747 38993
rect 3838 38757 4074 38993
rect 4165 38757 4401 38993
rect 4492 38757 4728 38993
rect 4819 38757 4967 38993
rect 4967 38757 5055 38993
rect 5146 38757 5382 38993
rect 5473 38757 5709 38993
rect 5800 38757 6036 38993
rect 6127 38757 6363 38993
rect 6454 38757 6690 38993
rect 6781 38757 7017 38993
rect 7108 38757 7344 38993
rect 7435 38757 7671 38993
rect 7762 38757 7998 38993
rect 8089 38757 8325 38993
rect 8415 38757 8651 38993
rect 8741 38757 8977 38993
rect 9067 38757 9303 38993
rect 9393 38757 9629 38993
rect 9719 38757 9955 38993
rect 10045 38757 10281 38993
rect 10371 38757 10607 38993
rect 10697 38757 10933 38993
rect 11023 38757 11259 38993
rect 11349 38757 11585 38993
rect 11675 38757 11911 38993
rect 12001 38757 12237 38993
rect 12327 38757 12563 38993
rect 12653 38757 12889 38993
rect 12979 38757 13215 38993
rect 13305 38757 13541 38993
rect 13631 38757 13867 38993
rect 13957 38757 14193 38993
rect 14283 38757 14519 38993
rect 14609 38757 14845 38993
rect 241 38433 477 38669
rect 568 38433 804 38669
rect 895 38433 1131 38669
rect 1222 38433 1458 38669
rect 1549 38433 1785 38669
rect 1876 38433 2112 38669
rect 2203 38433 2439 38669
rect 2530 38433 2766 38669
rect 2857 38433 3093 38669
rect 3184 38433 3420 38669
rect 3511 38433 3747 38669
rect 3838 38433 4074 38669
rect 4165 38433 4401 38669
rect 4492 38433 4728 38669
rect 4819 38433 4967 38669
rect 4967 38433 5055 38669
rect 5146 38433 5382 38669
rect 5473 38433 5709 38669
rect 5800 38433 6036 38669
rect 6127 38433 6363 38669
rect 6454 38433 6690 38669
rect 6781 38433 7017 38669
rect 7108 38433 7344 38669
rect 7435 38433 7671 38669
rect 7762 38433 7998 38669
rect 8089 38433 8325 38669
rect 8415 38433 8651 38669
rect 8741 38433 8977 38669
rect 9067 38433 9303 38669
rect 9393 38433 9629 38669
rect 9719 38433 9955 38669
rect 10045 38433 10281 38669
rect 10371 38433 10607 38669
rect 10697 38433 10933 38669
rect 11023 38433 11259 38669
rect 11349 38433 11585 38669
rect 11675 38433 11911 38669
rect 12001 38433 12237 38669
rect 12327 38433 12563 38669
rect 12653 38433 12889 38669
rect 12979 38433 13215 38669
rect 13305 38433 13541 38669
rect 13631 38433 13867 38669
rect 13957 38433 14193 38669
rect 14283 38433 14519 38669
rect 14609 38433 14845 38669
rect 241 38109 477 38345
rect 568 38109 804 38345
rect 895 38109 1131 38345
rect 1222 38109 1458 38345
rect 1549 38109 1785 38345
rect 1876 38109 2112 38345
rect 2203 38109 2439 38345
rect 2530 38109 2766 38345
rect 2857 38109 3093 38345
rect 3184 38109 3420 38345
rect 3511 38109 3747 38345
rect 3838 38109 4074 38345
rect 4165 38109 4401 38345
rect 4492 38109 4728 38345
rect 4819 38109 4967 38345
rect 4967 38109 5055 38345
rect 5146 38109 5382 38345
rect 5473 38109 5709 38345
rect 5800 38109 6036 38345
rect 6127 38109 6363 38345
rect 6454 38109 6690 38345
rect 6781 38109 7017 38345
rect 7108 38109 7344 38345
rect 7435 38109 7671 38345
rect 7762 38109 7998 38345
rect 8089 38109 8325 38345
rect 8415 38109 8651 38345
rect 8741 38109 8977 38345
rect 9067 38109 9303 38345
rect 9393 38109 9629 38345
rect 9719 38109 9955 38345
rect 10045 38109 10281 38345
rect 10371 38109 10607 38345
rect 10697 38109 10933 38345
rect 11023 38109 11259 38345
rect 11349 38109 11585 38345
rect 11675 38109 11911 38345
rect 12001 38109 12237 38345
rect 12327 38109 12563 38345
rect 12653 38109 12889 38345
rect 12979 38109 13215 38345
rect 13305 38109 13541 38345
rect 13631 38109 13867 38345
rect 13957 38109 14193 38345
rect 14283 38109 14519 38345
rect 14609 38109 14845 38345
rect 241 37785 477 38021
rect 568 37785 804 38021
rect 895 37785 1131 38021
rect 1222 37785 1458 38021
rect 1549 37785 1785 38021
rect 1876 37785 2112 38021
rect 2203 37785 2439 38021
rect 2530 37785 2766 38021
rect 2857 37785 3093 38021
rect 3184 37785 3420 38021
rect 3511 37785 3747 38021
rect 3838 37785 4074 38021
rect 4165 37785 4401 38021
rect 4492 37785 4728 38021
rect 4819 37785 4967 38021
rect 4967 37785 5055 38021
rect 5146 37785 5382 38021
rect 5473 37785 5709 38021
rect 5800 37785 6036 38021
rect 6127 37785 6363 38021
rect 6454 37785 6690 38021
rect 6781 37785 7017 38021
rect 7108 37785 7344 38021
rect 7435 37785 7671 38021
rect 7762 37785 7998 38021
rect 8089 37785 8325 38021
rect 8415 37785 8651 38021
rect 8741 37785 8977 38021
rect 9067 37785 9303 38021
rect 9393 37785 9629 38021
rect 9719 37785 9955 38021
rect 10045 37785 10281 38021
rect 10371 37785 10607 38021
rect 10697 37785 10933 38021
rect 11023 37785 11259 38021
rect 11349 37785 11585 38021
rect 11675 37785 11911 38021
rect 12001 37785 12237 38021
rect 12327 37785 12563 38021
rect 12653 37785 12889 38021
rect 12979 37785 13215 38021
rect 13305 37785 13541 38021
rect 13631 37785 13867 38021
rect 13957 37785 14193 38021
rect 14283 37785 14519 38021
rect 14609 37785 14845 38021
rect 241 37461 477 37697
rect 568 37461 804 37697
rect 895 37461 1131 37697
rect 1222 37461 1458 37697
rect 1549 37461 1785 37697
rect 1876 37461 2112 37697
rect 2203 37461 2439 37697
rect 2530 37461 2766 37697
rect 2857 37461 3093 37697
rect 3184 37461 3420 37697
rect 3511 37461 3747 37697
rect 3838 37461 4074 37697
rect 4165 37461 4401 37697
rect 4492 37461 4728 37697
rect 4819 37461 4967 37697
rect 4967 37461 5055 37697
rect 5146 37461 5382 37697
rect 5473 37461 5709 37697
rect 5800 37461 6036 37697
rect 6127 37461 6363 37697
rect 6454 37461 6690 37697
rect 6781 37461 7017 37697
rect 7108 37461 7344 37697
rect 7435 37461 7671 37697
rect 7762 37461 7998 37697
rect 8089 37461 8325 37697
rect 8415 37461 8651 37697
rect 8741 37461 8977 37697
rect 9067 37461 9303 37697
rect 9393 37461 9629 37697
rect 9719 37461 9955 37697
rect 10045 37461 10281 37697
rect 10371 37461 10607 37697
rect 10697 37461 10933 37697
rect 11023 37461 11259 37697
rect 11349 37461 11585 37697
rect 11675 37461 11911 37697
rect 12001 37461 12237 37697
rect 12327 37461 12563 37697
rect 12653 37461 12889 37697
rect 12979 37461 13215 37697
rect 13305 37461 13541 37697
rect 13631 37461 13867 37697
rect 13957 37461 14193 37697
rect 14283 37461 14519 37697
rect 14609 37461 14845 37697
rect 241 37137 477 37373
rect 568 37137 804 37373
rect 895 37198 1131 37373
rect 1222 37198 1458 37373
rect 1549 37198 1785 37373
rect 1876 37198 2112 37373
rect 895 37137 959 37198
rect 959 37137 1131 37198
rect 1222 37137 1458 37198
rect 1549 37137 1785 37198
rect 1876 37137 2112 37198
rect 2203 37137 2439 37373
rect 2530 37137 2766 37373
rect 2857 37137 3093 37373
rect 3184 37137 3420 37373
rect 3511 37137 3747 37373
rect 3838 37137 4074 37373
rect 4165 37137 4401 37373
rect 4492 37137 4728 37373
rect 4819 37137 4967 37373
rect 4967 37137 5055 37373
rect 5146 37137 5382 37373
rect 5473 37137 5709 37373
rect 5800 37137 6036 37373
rect 6127 37137 6363 37373
rect 6454 37137 6690 37373
rect 6781 37137 7017 37373
rect 7108 37137 7344 37373
rect 7435 37137 7671 37373
rect 7762 37137 7998 37373
rect 8089 37137 8325 37373
rect 8415 37137 8651 37373
rect 8741 37137 8977 37373
rect 9067 37137 9303 37373
rect 9393 37137 9629 37373
rect 9719 37137 9955 37373
rect 10045 37137 10281 37373
rect 10371 37137 10607 37373
rect 10697 37137 10933 37373
rect 11023 37137 11259 37373
rect 11349 37137 11585 37373
rect 11675 37137 11911 37373
rect 12001 37137 12237 37373
rect 12327 37137 12563 37373
rect 12653 37195 12889 37373
rect 12979 37195 13215 37373
rect 13305 37195 13541 37373
rect 13631 37195 13867 37373
rect 13957 37195 14193 37373
rect 12653 37137 12823 37195
rect 12823 37137 12889 37195
rect 12979 37137 13215 37195
rect 13305 37137 13541 37195
rect 13631 37137 13867 37195
rect 13957 37137 14007 37195
rect 14007 37137 14193 37195
rect 14283 37137 14519 37373
rect 14609 37137 14845 37373
rect 241 36813 477 37049
rect 568 36813 804 37049
rect 895 36813 959 37049
rect 959 36813 1131 37049
rect 1222 36813 1458 37049
rect 1549 36813 1785 37049
rect 1876 36813 2112 37049
rect 2203 36813 2439 37049
rect 2530 36813 2766 37049
rect 2857 36813 3093 37049
rect 3184 36813 3420 37049
rect 3511 36813 3747 37049
rect 3838 36813 4074 37049
rect 4165 36813 4401 37049
rect 4492 36813 4728 37049
rect 4819 36813 4967 37049
rect 4967 36813 5055 37049
rect 5146 36813 5382 37049
rect 5473 36813 5709 37049
rect 5800 36813 6036 37049
rect 6127 36813 6363 37049
rect 6454 36813 6690 37049
rect 6781 36813 7017 37049
rect 7108 36813 7344 37049
rect 7435 36813 7671 37049
rect 7762 36813 7998 37049
rect 8089 36813 8325 37049
rect 8415 36813 8651 37049
rect 8741 36813 8977 37049
rect 9067 36813 9303 37049
rect 9393 36813 9629 37049
rect 9719 36813 9955 37049
rect 10045 36813 10281 37049
rect 10371 36813 10607 37049
rect 10697 36813 10933 37049
rect 11023 36813 11259 37049
rect 11349 36813 11585 37049
rect 11675 36813 11911 37049
rect 12001 36813 12237 37049
rect 12327 36813 12563 37049
rect 12653 36813 12823 37049
rect 12823 36813 12889 37049
rect 12979 36813 13215 37049
rect 13305 36813 13541 37049
rect 13631 36813 13867 37049
rect 13957 36813 14007 37049
rect 14007 36813 14193 37049
rect 14283 36813 14519 37049
rect 14609 36813 14845 37049
rect 241 36489 477 36725
rect 568 36489 804 36725
rect 895 36494 959 36725
rect 959 36494 1131 36725
rect 1222 36494 1458 36725
rect 1549 36494 1785 36725
rect 1876 36494 2112 36725
rect 895 36489 1131 36494
rect 1222 36489 1458 36494
rect 1549 36489 1785 36494
rect 1876 36489 2112 36494
rect 2203 36489 2439 36725
rect 2530 36489 2766 36725
rect 2857 36489 3093 36725
rect 3184 36489 3420 36725
rect 3511 36489 3747 36725
rect 3838 36489 4074 36725
rect 4165 36489 4401 36725
rect 4492 36489 4728 36725
rect 4819 36489 4967 36725
rect 4967 36489 5055 36725
rect 5146 36489 5382 36725
rect 5473 36489 5709 36725
rect 5800 36489 6036 36725
rect 6127 36489 6363 36725
rect 6454 36489 6690 36725
rect 6781 36489 7017 36725
rect 7108 36489 7344 36725
rect 7435 36489 7671 36725
rect 7762 36489 7998 36725
rect 8089 36489 8325 36725
rect 8415 36489 8651 36725
rect 8741 36489 8977 36725
rect 9067 36489 9303 36725
rect 9393 36489 9629 36725
rect 9719 36489 9955 36725
rect 10045 36489 10281 36725
rect 10371 36489 10607 36725
rect 10697 36489 10933 36725
rect 11023 36489 11259 36725
rect 11349 36489 11585 36725
rect 11675 36489 11911 36725
rect 12001 36489 12237 36725
rect 12327 36489 12563 36725
rect 12653 36491 12823 36725
rect 12823 36491 12889 36725
rect 12979 36491 13215 36725
rect 13305 36491 13541 36725
rect 13631 36491 13867 36725
rect 13957 36491 14007 36725
rect 14007 36491 14193 36725
rect 12653 36489 12889 36491
rect 12979 36489 13215 36491
rect 13305 36489 13541 36491
rect 13631 36489 13867 36491
rect 13957 36489 14193 36491
rect 14283 36489 14519 36725
rect 14609 36489 14845 36725
rect 241 36165 477 36401
rect 568 36165 804 36401
rect 895 36165 1131 36401
rect 1222 36165 1458 36401
rect 1549 36165 1785 36401
rect 1876 36165 2112 36401
rect 2203 36165 2439 36401
rect 2530 36165 2766 36401
rect 2857 36165 3093 36401
rect 3184 36165 3420 36401
rect 3511 36165 3747 36401
rect 3838 36165 4074 36401
rect 4165 36165 4401 36401
rect 4492 36165 4728 36401
rect 4819 36165 4967 36401
rect 4967 36165 5055 36401
rect 5146 36165 5382 36401
rect 5473 36165 5709 36401
rect 5800 36165 6036 36401
rect 6127 36165 6363 36401
rect 6454 36165 6690 36401
rect 6781 36165 7017 36401
rect 7108 36165 7344 36401
rect 7435 36165 7671 36401
rect 7762 36165 7998 36401
rect 8089 36165 8325 36401
rect 8415 36165 8651 36401
rect 8741 36165 8977 36401
rect 9067 36165 9303 36401
rect 9393 36165 9629 36401
rect 9719 36165 9955 36401
rect 10045 36165 10281 36401
rect 10371 36165 10607 36401
rect 10697 36165 10933 36401
rect 11023 36165 11259 36401
rect 11349 36165 11585 36401
rect 11675 36165 11911 36401
rect 12001 36165 12237 36401
rect 12327 36165 12563 36401
rect 12653 36165 12889 36401
rect 12979 36165 13215 36401
rect 13305 36165 13541 36401
rect 13631 36165 13867 36401
rect 13957 36165 14193 36401
rect 14283 36165 14519 36401
rect 14609 36165 14845 36401
rect 241 35841 477 36077
rect 568 35841 804 36077
rect 895 35841 1131 36077
rect 1222 35841 1458 36077
rect 1549 35841 1785 36077
rect 1876 35841 2112 36077
rect 2203 35841 2439 36077
rect 2530 35841 2766 36077
rect 2857 35841 3093 36077
rect 3184 35841 3420 36077
rect 3511 35841 3747 36077
rect 3838 35841 4074 36077
rect 4165 35841 4401 36077
rect 4492 35841 4728 36077
rect 4819 35841 4967 36077
rect 4967 35841 5055 36077
rect 5146 35841 5382 36077
rect 5473 35841 5709 36077
rect 5800 35841 6036 36077
rect 6127 35841 6363 36077
rect 6454 35841 6690 36077
rect 6781 35841 7017 36077
rect 7108 35841 7344 36077
rect 7435 35841 7671 36077
rect 7762 35841 7998 36077
rect 8089 35841 8325 36077
rect 8415 35841 8651 36077
rect 8741 35841 8977 36077
rect 9067 35841 9303 36077
rect 9393 35841 9629 36077
rect 9719 35841 9955 36077
rect 10045 35841 10281 36077
rect 10371 35841 10607 36077
rect 10697 35841 10933 36077
rect 11023 35841 11259 36077
rect 11349 35841 11585 36077
rect 11675 35841 11911 36077
rect 12001 35841 12237 36077
rect 12327 35841 12563 36077
rect 12653 35841 12889 36077
rect 12979 35841 13215 36077
rect 13305 35841 13541 36077
rect 13631 35841 13867 36077
rect 13957 35841 14193 36077
rect 14283 35841 14519 36077
rect 14609 35841 14845 36077
rect 241 35517 477 35753
rect 568 35517 804 35753
rect 895 35517 1131 35753
rect 1222 35517 1458 35753
rect 1549 35517 1785 35753
rect 1876 35517 2112 35753
rect 2203 35517 2439 35753
rect 2530 35517 2766 35753
rect 2857 35517 3093 35753
rect 3184 35517 3420 35753
rect 3511 35517 3747 35753
rect 3838 35517 4074 35753
rect 4165 35517 4401 35753
rect 4492 35517 4728 35753
rect 4819 35517 4967 35753
rect 4967 35517 5055 35753
rect 5146 35517 5382 35753
rect 5473 35517 5709 35753
rect 5800 35517 6036 35753
rect 6127 35517 6363 35753
rect 6454 35517 6690 35753
rect 6781 35517 7017 35753
rect 7108 35517 7344 35753
rect 7435 35517 7671 35753
rect 7762 35517 7998 35753
rect 8089 35517 8325 35753
rect 8415 35517 8651 35753
rect 8741 35517 8977 35753
rect 9067 35517 9303 35753
rect 9393 35517 9629 35753
rect 9719 35517 9955 35753
rect 10045 35517 10281 35753
rect 10371 35517 10607 35753
rect 10697 35517 10933 35753
rect 11023 35517 11259 35753
rect 11349 35517 11585 35753
rect 11675 35517 11911 35753
rect 12001 35517 12237 35753
rect 12327 35517 12563 35753
rect 12653 35517 12889 35753
rect 12979 35517 13215 35753
rect 13305 35517 13541 35753
rect 13631 35517 13867 35753
rect 13957 35517 14193 35753
rect 14283 35517 14519 35753
rect 14609 35517 14845 35753
rect 241 35193 477 35429
rect 568 35193 804 35429
rect 895 35193 1131 35429
rect 1222 35193 1458 35429
rect 1549 35193 1785 35429
rect 1876 35193 2112 35429
rect 2203 35193 2439 35429
rect 2530 35193 2766 35429
rect 2857 35193 3093 35429
rect 3184 35193 3420 35429
rect 3511 35193 3747 35429
rect 3838 35193 4074 35429
rect 4165 35193 4401 35429
rect 4492 35193 4728 35429
rect 4819 35324 4967 35429
rect 4967 35324 5055 35429
rect 5146 35324 5382 35429
rect 5473 35324 5709 35429
rect 5800 35324 6036 35429
rect 6127 35324 6363 35429
rect 6454 35324 6690 35429
rect 6781 35324 7017 35429
rect 7108 35324 7344 35429
rect 7435 35324 7671 35429
rect 7762 35324 7998 35429
rect 8089 35324 8325 35429
rect 8415 35324 8651 35429
rect 8741 35324 8977 35429
rect 9067 35324 9303 35429
rect 9393 35324 9629 35429
rect 9719 35324 9955 35429
rect 4819 35193 5055 35324
rect 5146 35193 5382 35324
rect 5473 35193 5709 35324
rect 5800 35193 6036 35324
rect 6127 35193 6363 35324
rect 6454 35193 6690 35324
rect 6781 35193 7017 35324
rect 7108 35193 7344 35324
rect 7435 35193 7671 35324
rect 7762 35193 7998 35324
rect 8089 35193 8325 35324
rect 8415 35193 8651 35324
rect 8741 35193 8977 35324
rect 9067 35193 9303 35324
rect 9393 35193 9629 35324
rect 9719 35193 9955 35324
rect 10045 35193 10281 35429
rect 10371 35193 10607 35429
rect 10697 35193 10933 35429
rect 11023 35193 11259 35429
rect 11349 35193 11585 35429
rect 11675 35193 11911 35429
rect 12001 35193 12237 35429
rect 12327 35193 12563 35429
rect 12653 35193 12889 35429
rect 12979 35193 13215 35429
rect 13305 35193 13541 35429
rect 13631 35193 13867 35429
rect 13957 35193 14193 35429
rect 14283 35193 14519 35429
rect 14609 35193 14845 35429
rect 2268 34588 2504 34596
rect 2588 34588 2824 34596
rect 2908 34588 3144 34596
rect 2268 34360 2331 34588
rect 2331 34360 2504 34588
rect 2588 34360 2824 34588
rect 2908 34360 3035 34588
rect 3035 34360 3144 34588
rect 3228 34360 3464 34596
rect 3548 34360 3784 34596
rect 3868 34360 4104 34596
rect 4188 34360 4424 34596
rect 4508 34360 4744 34596
rect 4828 34360 5064 34596
rect 5148 34360 5384 34596
rect 5468 34360 5704 34596
rect 5788 34360 6024 34596
rect 6108 34360 6344 34596
rect 6428 34360 6664 34596
rect 6748 34360 6984 34596
rect 7068 34360 7304 34596
rect 7388 34360 7624 34596
rect 7708 34360 7944 34596
rect 8028 34360 8264 34596
rect 8348 34360 8584 34596
rect 8668 34360 8904 34596
rect 8988 34360 9224 34596
rect 9308 34360 9544 34596
rect 9628 34360 9864 34596
rect 9948 34360 10184 34596
rect 10268 34360 10504 34596
rect 10588 34360 10824 34596
rect 10908 34360 11144 34596
rect 11228 34360 11464 34596
rect 11548 34360 11784 34596
rect 11868 34587 12104 34596
rect 12188 34587 12424 34596
rect 12508 34587 12744 34596
rect 11868 34360 11961 34587
rect 11961 34360 12104 34587
rect 12188 34360 12424 34587
rect 12508 34360 12665 34587
rect 12665 34360 12744 34587
rect 1946 34052 2182 34288
rect 1626 33732 1862 33968
rect 12870 33998 13106 34234
rect 1306 33412 1542 33648
rect 983 33089 1219 33325
rect 13190 33678 13426 33914
rect 13510 33358 13746 33594
rect 983 32974 1219 33005
rect 983 32769 1035 32974
rect 1035 32769 1219 32974
rect 983 32449 1035 32685
rect 1035 32449 1219 32685
rect 983 32129 1035 32365
rect 1035 32129 1219 32365
rect 983 31809 1035 32045
rect 1035 31809 1219 32045
rect 983 31489 1035 31725
rect 1035 31489 1219 31725
rect 983 31169 1035 31405
rect 1035 31169 1219 31405
rect 983 30849 1035 31085
rect 1035 30849 1219 31085
rect 983 30529 1035 30765
rect 1035 30529 1219 30765
rect 983 30209 1035 30445
rect 1035 30209 1219 30445
rect 983 29889 1035 30125
rect 1035 29889 1219 30125
rect 983 29569 1035 29805
rect 1035 29569 1219 29805
rect 983 29249 1035 29485
rect 1035 29249 1219 29485
rect 983 28929 1035 29165
rect 1035 28929 1219 29165
rect 983 28609 1035 28845
rect 1035 28609 1219 28845
rect 983 28289 1035 28525
rect 1035 28289 1219 28525
rect 983 27969 1035 28205
rect 1035 27969 1219 28205
rect 983 27649 1035 27885
rect 1035 27649 1219 27885
rect 983 27329 1035 27565
rect 1035 27329 1219 27565
rect 983 27009 1035 27245
rect 1035 27009 1219 27245
rect 983 26689 1035 26925
rect 1035 26689 1219 26925
rect 983 26369 1035 26605
rect 1035 26369 1219 26605
rect 983 26049 1035 26285
rect 1035 26049 1219 26285
rect 983 25729 1035 25965
rect 1035 25729 1219 25965
rect 983 25409 1035 25645
rect 1035 25409 1219 25645
rect 983 25089 1035 25325
rect 1035 25089 1219 25325
rect 983 24769 1035 25005
rect 1035 24769 1219 25005
rect 983 24449 1035 24685
rect 1035 24449 1219 24685
rect 983 24129 1035 24365
rect 1035 24129 1219 24365
rect 983 23809 1035 24045
rect 1035 23809 1219 24045
rect 983 23489 1035 23725
rect 1035 23489 1219 23725
rect 983 23169 1035 23405
rect 1035 23169 1219 23405
rect 983 22849 1035 23085
rect 1035 22849 1219 23085
rect 983 22529 1035 22765
rect 1035 22529 1219 22765
rect 983 22209 1035 22445
rect 1035 22209 1219 22445
rect 983 21889 1035 22125
rect 1035 21889 1219 22125
rect 983 21569 1035 21805
rect 1035 21569 1219 21805
rect 983 21249 1035 21485
rect 1035 21249 1219 21485
rect 983 20929 1219 21165
rect 13779 32995 14015 33231
rect 13779 32866 14015 32911
rect 13779 32675 13965 32866
rect 13965 32675 14015 32866
rect 13779 32355 13965 32591
rect 13965 32355 14015 32591
rect 13779 32035 13965 32271
rect 13965 32035 14015 32271
rect 13779 31715 13965 31951
rect 13965 31715 14015 31951
rect 13779 31395 13965 31631
rect 13965 31395 14015 31631
rect 13779 31075 13965 31311
rect 13965 31075 14015 31311
rect 13779 30755 13965 30991
rect 13965 30755 14015 30991
rect 13779 30435 13965 30671
rect 13965 30435 14015 30671
rect 13779 30115 13965 30351
rect 13965 30115 14015 30351
rect 13779 29795 13965 30031
rect 13965 29795 14015 30031
rect 13779 29475 13965 29711
rect 13965 29475 14015 29711
rect 13779 29155 13965 29391
rect 13965 29155 14015 29391
rect 13779 28835 13965 29071
rect 13965 28835 14015 29071
rect 13779 28515 13965 28751
rect 13965 28515 14015 28751
rect 13779 28195 13965 28431
rect 13965 28195 14015 28431
rect 13779 27875 13965 28111
rect 13965 27875 14015 28111
rect 13779 27555 13965 27791
rect 13965 27555 14015 27791
rect 13779 27235 13965 27471
rect 13965 27235 14015 27471
rect 13779 26915 13965 27151
rect 13965 26915 14015 27151
rect 13779 26595 13965 26831
rect 13965 26595 14015 26831
rect 13779 26275 13965 26511
rect 13965 26275 14015 26511
rect 13779 25955 13965 26191
rect 13965 25955 14015 26191
rect 13779 25635 13965 25871
rect 13965 25635 14015 25871
rect 13779 25315 13965 25551
rect 13965 25315 14015 25551
rect 13779 24995 13965 25231
rect 13965 24995 14015 25231
rect 13779 24675 13965 24911
rect 13965 24675 14015 24911
rect 13779 24355 13965 24591
rect 13965 24355 14015 24591
rect 13779 24035 13965 24271
rect 13965 24035 14015 24271
rect 13779 23715 13965 23951
rect 13965 23715 14015 23951
rect 13779 23395 13965 23631
rect 13965 23395 14015 23631
rect 13779 23075 13965 23311
rect 13965 23075 14015 23311
rect 13779 22755 13965 22991
rect 13965 22755 14015 22991
rect 13779 22435 13965 22671
rect 13965 22435 14015 22671
rect 13779 22115 13965 22351
rect 13965 22115 14015 22351
rect 13779 21795 13965 22031
rect 13965 21795 14015 22031
rect 13779 21475 13965 21711
rect 13965 21475 14015 21711
rect 13779 21155 13965 21391
rect 13965 21155 14015 21391
rect 1252 20566 1488 20802
rect 1572 20246 1808 20482
rect 13779 20835 14015 21071
rect 13456 20512 13692 20748
rect 1892 19926 2128 20162
rect 13136 20192 13372 20428
rect 12816 19872 13052 20108
rect 2254 19576 2308 19800
rect 2308 19576 2490 19800
rect 2574 19576 2810 19800
rect 2894 19576 3130 19800
rect 3214 19576 3450 19800
rect 3534 19576 3770 19800
rect 3854 19576 4090 19800
rect 4174 19576 4410 19800
rect 4494 19576 4730 19800
rect 4814 19576 5050 19800
rect 5134 19576 5370 19800
rect 5454 19576 5690 19800
rect 5774 19576 6010 19800
rect 6094 19576 6330 19800
rect 6414 19576 6650 19800
rect 6734 19576 6970 19800
rect 7054 19576 7290 19800
rect 7374 19576 7610 19800
rect 7694 19576 7930 19800
rect 8014 19576 8250 19800
rect 8334 19576 8570 19800
rect 8654 19576 8890 19800
rect 8974 19576 9210 19800
rect 9294 19576 9530 19800
rect 9614 19576 9850 19800
rect 9934 19576 10170 19800
rect 10254 19576 10490 19800
rect 10574 19576 10810 19800
rect 10894 19576 11130 19800
rect 11214 19576 11450 19800
rect 11534 19576 11770 19800
rect 11854 19576 12090 19800
rect 12174 19576 12410 19800
rect 12494 19576 12692 19800
rect 12692 19576 12730 19800
rect 2254 19564 2490 19576
rect 2574 19564 2810 19576
rect 2894 19564 3130 19576
rect 3214 19564 3450 19576
rect 3534 19564 3770 19576
rect 3854 19564 4090 19576
rect 4174 19564 4410 19576
rect 4494 19564 4730 19576
rect 4814 19564 5050 19576
rect 5134 19564 5370 19576
rect 5454 19564 5690 19576
rect 5774 19564 6010 19576
rect 6094 19564 6330 19576
rect 6414 19564 6650 19576
rect 6734 19564 6970 19576
rect 7054 19564 7290 19576
rect 7374 19564 7610 19576
rect 7694 19564 7930 19576
rect 8014 19564 8250 19576
rect 8334 19564 8570 19576
rect 8654 19564 8890 19576
rect 8974 19564 9210 19576
rect 9294 19564 9530 19576
rect 9614 19564 9850 19576
rect 9934 19564 10170 19576
rect 10254 19564 10490 19576
rect 10574 19564 10810 19576
rect 10894 19564 11130 19576
rect 11214 19564 11450 19576
rect 11534 19564 11770 19576
rect 11854 19564 12090 19576
rect 12174 19564 12410 19576
rect 12494 19564 12730 19576
rect 143 18736 379 18972
rect 465 18736 701 18972
rect 787 18736 1023 18972
rect 1109 18736 1345 18972
rect 1431 18736 1667 18972
rect 1753 18736 1989 18972
rect 2075 18736 2311 18972
rect 2397 18736 2633 18972
rect 2719 18908 2955 18972
rect 3041 18908 3277 18972
rect 3363 18908 3599 18972
rect 3685 18908 3921 18972
rect 4007 18908 4243 18972
rect 4329 18908 4565 18972
rect 4651 18908 4887 18972
rect 4973 18908 5209 18972
rect 2719 18736 2930 18908
rect 2930 18736 2955 18908
rect 3041 18736 3277 18908
rect 3363 18736 3599 18908
rect 3685 18736 3921 18908
rect 4007 18736 4243 18908
rect 4329 18736 4565 18908
rect 4651 18736 4887 18908
rect 4973 18736 5209 18908
rect 5295 18736 5531 18972
rect 143 18400 379 18636
rect 465 18400 701 18636
rect 787 18400 1023 18636
rect 1109 18400 1345 18636
rect 1431 18400 1667 18636
rect 1753 18400 1989 18636
rect 2075 18400 2311 18636
rect 2397 18400 2633 18636
rect 2719 18400 2930 18636
rect 2930 18400 2955 18636
rect 3041 18400 3277 18636
rect 3363 18400 3599 18636
rect 3685 18400 3921 18636
rect 4007 18400 4243 18636
rect 4329 18400 4565 18636
rect 4651 18400 4887 18636
rect 4973 18400 5209 18636
rect 5295 18400 5531 18636
rect 143 18064 379 18300
rect 465 18064 701 18300
rect 787 18064 1023 18300
rect 1109 18064 1345 18300
rect 1431 18064 1667 18300
rect 1753 18064 1989 18300
rect 2075 18064 2311 18300
rect 2397 18064 2633 18300
rect 2719 18064 2930 18300
rect 2930 18064 2955 18300
rect 3041 18064 3277 18300
rect 3363 18064 3599 18300
rect 3685 18064 3921 18300
rect 4007 18064 4243 18300
rect 4329 18064 4565 18300
rect 4651 18064 4887 18300
rect 4973 18064 5209 18300
rect 5295 18064 5531 18300
rect 143 17728 379 17964
rect 465 17728 701 17964
rect 787 17728 1023 17964
rect 1109 17728 1345 17964
rect 1431 17728 1667 17964
rect 1753 17728 1989 17964
rect 2075 17728 2311 17964
rect 2397 17728 2633 17964
rect 2719 17728 2930 17964
rect 2930 17728 2955 17964
rect 3041 17728 3277 17964
rect 3363 17728 3599 17964
rect 3685 17728 3921 17964
rect 4007 17728 4243 17964
rect 4329 17728 4565 17964
rect 4651 17728 4887 17964
rect 4973 17728 5209 17964
rect 5295 17728 5531 17964
rect 143 17392 379 17628
rect 465 17392 701 17628
rect 787 17392 1023 17628
rect 1109 17392 1345 17628
rect 1431 17392 1667 17628
rect 1753 17392 1989 17628
rect 2075 17392 2311 17628
rect 2397 17392 2633 17628
rect 2719 17392 2930 17628
rect 2930 17392 2955 17628
rect 3041 17392 3277 17628
rect 3363 17392 3599 17628
rect 3685 17392 3921 17628
rect 4007 17392 4243 17628
rect 4329 17392 4565 17628
rect 4651 17392 4887 17628
rect 4973 17392 5209 17628
rect 5295 17392 5531 17628
rect 143 17056 379 17292
rect 465 17056 701 17292
rect 787 17056 1023 17292
rect 1109 17056 1345 17292
rect 1431 17056 1667 17292
rect 1753 17056 1989 17292
rect 2075 17056 2311 17292
rect 2397 17056 2633 17292
rect 2719 17056 2955 17292
rect 3041 17231 3277 17292
rect 3363 17231 3599 17292
rect 3685 17231 3921 17292
rect 4007 17231 4243 17292
rect 4329 17231 4565 17292
rect 4651 17231 4887 17292
rect 4973 17231 5209 17292
rect 3041 17087 3091 17231
rect 3091 17087 3277 17231
rect 3363 17087 3599 17231
rect 3685 17087 3921 17231
rect 4007 17087 4243 17231
rect 4329 17087 4565 17231
rect 4651 17087 4887 17231
rect 4973 17087 5209 17231
rect 3041 17056 3277 17087
rect 3363 17056 3599 17087
rect 3685 17056 3921 17087
rect 4007 17056 4243 17087
rect 4329 17056 4565 17087
rect 4651 17056 4887 17087
rect 4973 17056 5209 17087
rect 5295 17056 5531 17292
rect 143 16720 379 16956
rect 465 16720 701 16956
rect 787 16720 1023 16956
rect 1109 16720 1345 16956
rect 1431 16720 1667 16956
rect 1753 16720 1989 16956
rect 2075 16720 2311 16956
rect 2397 16720 2633 16956
rect 2719 16720 2955 16956
rect 3041 16720 3277 16956
rect 3363 16720 3599 16956
rect 3685 16720 3921 16956
rect 4007 16720 4243 16956
rect 4329 16720 4565 16956
rect 4651 16720 4887 16956
rect 4973 16720 5209 16956
rect 5295 16720 5531 16956
rect 143 16384 379 16620
rect 465 16384 701 16620
rect 787 16384 1023 16620
rect 1109 16384 1345 16620
rect 1431 16384 1667 16620
rect 1753 16384 1989 16620
rect 2075 16384 2311 16620
rect 2397 16384 2633 16620
rect 2719 16384 2955 16620
rect 3041 16384 3277 16620
rect 3363 16384 3599 16620
rect 3685 16384 3921 16620
rect 4007 16384 4243 16620
rect 4329 16384 4565 16620
rect 4651 16384 4887 16620
rect 4973 16384 5209 16620
rect 5295 16384 5531 16620
rect 143 16048 379 16284
rect 465 16048 701 16284
rect 787 16048 1023 16284
rect 1109 16048 1345 16284
rect 1431 16048 1667 16284
rect 1753 16048 1989 16284
rect 2075 16048 2311 16284
rect 2397 16048 2633 16284
rect 2719 16048 2955 16284
rect 3041 16048 3277 16284
rect 3363 16048 3599 16284
rect 3685 16048 3921 16284
rect 4007 16048 4243 16284
rect 4329 16048 4565 16284
rect 4651 16048 4887 16284
rect 4973 16048 5209 16284
rect 5295 16048 5531 16284
rect 143 15712 379 15948
rect 465 15712 701 15948
rect 787 15712 1023 15948
rect 1109 15712 1345 15948
rect 1431 15712 1667 15948
rect 1753 15712 1989 15948
rect 2075 15712 2311 15948
rect 2397 15712 2633 15948
rect 2719 15712 2955 15948
rect 3041 15712 3277 15948
rect 3363 15712 3599 15948
rect 3685 15712 3921 15948
rect 4007 15712 4243 15948
rect 4329 15712 4565 15948
rect 4651 15712 4887 15948
rect 4973 15712 5209 15948
rect 5295 15712 5531 15948
rect 143 15376 379 15612
rect 465 15376 701 15612
rect 787 15376 1023 15612
rect 1109 15376 1345 15612
rect 1431 15376 1667 15612
rect 1753 15376 1989 15612
rect 2075 15376 2311 15612
rect 2397 15376 2633 15612
rect 2719 15376 2955 15612
rect 3041 15376 3277 15612
rect 3363 15376 3599 15612
rect 3685 15376 3921 15612
rect 4007 15376 4243 15612
rect 4329 15376 4565 15612
rect 4651 15376 4887 15612
rect 4973 15376 5209 15612
rect 5295 15376 5531 15612
rect 143 15040 379 15276
rect 465 15040 701 15276
rect 787 15040 1023 15276
rect 1109 15040 1345 15276
rect 1431 15040 1667 15276
rect 1753 15040 1989 15276
rect 2075 15040 2311 15276
rect 2397 15040 2633 15276
rect 2719 15040 2955 15276
rect 3041 15040 3277 15276
rect 3363 15040 3599 15276
rect 3685 15040 3921 15276
rect 4007 15040 4243 15276
rect 4329 15040 4565 15276
rect 4651 15040 4887 15276
rect 4973 15040 5209 15276
rect 5295 15040 5531 15276
rect 143 14704 379 14940
rect 465 14704 701 14940
rect 787 14718 1023 14940
rect 1109 14718 1345 14940
rect 1431 14718 1667 14940
rect 1753 14718 1989 14940
rect 787 14704 918 14718
rect 918 14704 1023 14718
rect 1109 14704 1345 14718
rect 1431 14704 1667 14718
rect 1753 14704 1989 14718
rect 2075 14704 2311 14940
rect 2397 14704 2633 14940
rect 2719 14704 2955 14940
rect 3041 14704 3277 14940
rect 3363 14704 3599 14940
rect 3685 14704 3921 14940
rect 4007 14704 4243 14940
rect 4329 14704 4565 14940
rect 4651 14704 4887 14940
rect 4973 14704 5209 14940
rect 5295 14704 5531 14940
rect 143 14368 379 14604
rect 465 14368 701 14604
rect 787 14368 918 14604
rect 918 14368 1023 14604
rect 1109 14368 1345 14604
rect 1431 14368 1667 14604
rect 1753 14368 1989 14604
rect 2075 14368 2311 14604
rect 2397 14368 2633 14604
rect 2719 14368 2955 14604
rect 3041 14368 3277 14604
rect 3363 14368 3599 14604
rect 3685 14368 3921 14604
rect 4007 14368 4243 14604
rect 4329 14368 4565 14604
rect 4651 14368 4887 14604
rect 4973 14368 5209 14604
rect 5295 14368 5531 14604
rect 143 14032 379 14268
rect 465 14032 701 14268
rect 787 14032 1023 14268
rect 1109 14032 1345 14268
rect 1431 14032 1667 14268
rect 1753 14032 1989 14268
rect 2075 14032 2311 14268
rect 2397 14032 2633 14268
rect 2719 14032 2955 14268
rect 3041 14032 3277 14268
rect 3363 14032 3599 14268
rect 3685 14032 3921 14268
rect 4007 14032 4243 14268
rect 4329 14032 4565 14268
rect 4651 14032 4887 14268
rect 4973 14032 5209 14268
rect 5295 14032 5531 14268
rect 9469 18736 9705 18972
rect 9790 18908 10026 18972
rect 10111 18908 10347 18972
rect 10432 18908 10668 18972
rect 10753 18908 10989 18972
rect 11074 18908 11310 18972
rect 11395 18908 11631 18972
rect 11716 18908 11952 18972
rect 9790 18736 10026 18908
rect 10111 18736 10347 18908
rect 10432 18736 10668 18908
rect 10753 18736 10989 18908
rect 11074 18736 11310 18908
rect 11395 18736 11631 18908
rect 11716 18736 11952 18908
rect 12037 18736 12273 18972
rect 12358 18736 12594 18972
rect 12679 18736 12915 18972
rect 13000 18736 13236 18972
rect 13321 18736 13557 18972
rect 13642 18736 13878 18972
rect 13963 18736 14199 18972
rect 14284 18736 14520 18972
rect 14605 18736 14841 18972
rect 9469 18400 9705 18636
rect 9790 18400 10026 18636
rect 10111 18400 10347 18636
rect 10432 18400 10668 18636
rect 10753 18400 10989 18636
rect 11074 18400 11310 18636
rect 11395 18400 11631 18636
rect 11716 18400 11952 18636
rect 12037 18400 12273 18636
rect 12358 18400 12594 18636
rect 12679 18400 12915 18636
rect 13000 18400 13236 18636
rect 13321 18400 13557 18636
rect 13642 18400 13878 18636
rect 13963 18400 14199 18636
rect 14284 18400 14520 18636
rect 14605 18400 14841 18636
rect 9469 18064 9705 18300
rect 9790 18064 10026 18300
rect 10111 18064 10347 18300
rect 10432 18064 10668 18300
rect 10753 18064 10989 18300
rect 11074 18064 11310 18300
rect 11395 18064 11631 18300
rect 11716 18064 11952 18300
rect 12037 18064 12273 18300
rect 12358 18064 12594 18300
rect 12679 18064 12915 18300
rect 13000 18064 13236 18300
rect 13321 18064 13557 18300
rect 13642 18064 13878 18300
rect 13963 18064 14199 18300
rect 14284 18064 14520 18300
rect 14605 18064 14841 18300
rect 9469 17728 9705 17964
rect 9790 17728 10026 17964
rect 10111 17728 10347 17964
rect 10432 17728 10668 17964
rect 10753 17728 10989 17964
rect 11074 17728 11310 17964
rect 11395 17728 11631 17964
rect 11716 17728 11952 17964
rect 12037 17728 12273 17964
rect 12358 17728 12594 17964
rect 12679 17728 12915 17964
rect 13000 17728 13236 17964
rect 13321 17728 13557 17964
rect 13642 17728 13878 17964
rect 13963 17728 14199 17964
rect 14284 17728 14520 17964
rect 14605 17728 14841 17964
rect 9469 17392 9705 17628
rect 9790 17392 10026 17628
rect 10111 17392 10347 17628
rect 10432 17392 10668 17628
rect 10753 17392 10989 17628
rect 11074 17392 11310 17628
rect 11395 17392 11631 17628
rect 11716 17392 11952 17628
rect 12037 17392 12273 17628
rect 12358 17392 12594 17628
rect 12679 17392 12915 17628
rect 13000 17392 13236 17628
rect 13321 17392 13557 17628
rect 13642 17392 13878 17628
rect 13963 17392 14199 17628
rect 14284 17392 14520 17628
rect 14605 17392 14841 17628
rect 9469 17056 9705 17292
rect 9790 17231 10026 17292
rect 10111 17231 10347 17292
rect 10432 17231 10668 17292
rect 10753 17231 10989 17292
rect 11074 17231 11310 17292
rect 11395 17231 11631 17292
rect 11716 17231 11952 17292
rect 9790 17087 10026 17231
rect 10111 17087 10347 17231
rect 10432 17087 10668 17231
rect 10753 17087 10989 17231
rect 11074 17087 11310 17231
rect 11395 17087 11631 17231
rect 11716 17087 11871 17231
rect 11871 17087 11952 17231
rect 9790 17056 10026 17087
rect 10111 17056 10347 17087
rect 10432 17056 10668 17087
rect 10753 17056 10989 17087
rect 11074 17056 11310 17087
rect 11395 17056 11631 17087
rect 11716 17056 11952 17087
rect 12037 17056 12273 17292
rect 12358 17056 12594 17292
rect 12679 17056 12915 17292
rect 13000 17056 13236 17292
rect 13321 17056 13557 17292
rect 13642 17056 13878 17292
rect 13963 17056 14199 17292
rect 14284 17056 14520 17292
rect 14605 17056 14841 17292
rect 9469 16720 9705 16956
rect 9790 16720 10026 16956
rect 10111 16720 10347 16956
rect 10432 16720 10668 16956
rect 10753 16720 10989 16956
rect 11074 16720 11310 16956
rect 11395 16720 11631 16956
rect 11716 16720 11952 16956
rect 12037 16720 12273 16956
rect 12358 16720 12594 16956
rect 12679 16720 12915 16956
rect 13000 16720 13236 16956
rect 13321 16720 13557 16956
rect 13642 16720 13878 16956
rect 13963 16720 14199 16956
rect 14284 16720 14520 16956
rect 14605 16720 14841 16956
rect 9469 16384 9705 16620
rect 9790 16384 10026 16620
rect 10111 16384 10347 16620
rect 10432 16384 10668 16620
rect 10753 16384 10989 16620
rect 11074 16384 11310 16620
rect 11395 16384 11631 16620
rect 11716 16384 11952 16620
rect 12037 16384 12273 16620
rect 12358 16384 12594 16620
rect 12679 16384 12915 16620
rect 13000 16384 13236 16620
rect 13321 16384 13557 16620
rect 13642 16384 13878 16620
rect 13963 16384 14199 16620
rect 14284 16384 14520 16620
rect 14605 16384 14841 16620
rect 9469 16048 9705 16284
rect 9790 16048 10026 16284
rect 10111 16048 10347 16284
rect 10432 16048 10668 16284
rect 10753 16048 10989 16284
rect 11074 16048 11310 16284
rect 11395 16048 11631 16284
rect 11716 16048 11952 16284
rect 12037 16048 12273 16284
rect 12358 16048 12594 16284
rect 12679 16048 12915 16284
rect 13000 16048 13236 16284
rect 13321 16048 13557 16284
rect 13642 16048 13878 16284
rect 13963 16048 14199 16284
rect 14284 16048 14520 16284
rect 14605 16048 14841 16284
rect 9469 15712 9705 15948
rect 9790 15712 10026 15948
rect 10111 15712 10347 15948
rect 10432 15712 10668 15948
rect 10753 15712 10989 15948
rect 11074 15712 11310 15948
rect 11395 15712 11631 15948
rect 11716 15712 11952 15948
rect 12037 15712 12273 15948
rect 12358 15712 12594 15948
rect 12679 15712 12915 15948
rect 13000 15712 13236 15948
rect 13321 15712 13557 15948
rect 13642 15712 13878 15948
rect 13963 15712 14199 15948
rect 14284 15712 14520 15948
rect 14605 15712 14841 15948
rect 9469 15376 9705 15612
rect 9790 15376 10026 15612
rect 10111 15376 10347 15612
rect 10432 15376 10668 15612
rect 10753 15376 10989 15612
rect 11074 15376 11310 15612
rect 11395 15376 11631 15612
rect 11716 15376 11952 15612
rect 12037 15376 12273 15612
rect 12358 15376 12594 15612
rect 12679 15376 12915 15612
rect 13000 15376 13236 15612
rect 13321 15376 13557 15612
rect 13642 15376 13878 15612
rect 13963 15376 14199 15612
rect 14284 15376 14520 15612
rect 14605 15376 14841 15612
rect 9469 15040 9705 15276
rect 9790 15040 10026 15276
rect 10111 15040 10347 15276
rect 10432 15040 10668 15276
rect 10753 15040 10989 15276
rect 11074 15040 11310 15276
rect 11395 15040 11631 15276
rect 11716 15040 11952 15276
rect 12037 15040 12273 15276
rect 12358 15040 12594 15276
rect 12679 15040 12915 15276
rect 13000 15040 13236 15276
rect 13321 15040 13557 15276
rect 13642 15040 13878 15276
rect 13963 15040 14199 15276
rect 14284 15040 14520 15276
rect 14605 15040 14841 15276
rect 9469 14704 9705 14940
rect 9790 14704 10026 14940
rect 10111 14704 10347 14940
rect 10432 14704 10668 14940
rect 10753 14704 10989 14940
rect 11074 14704 11310 14940
rect 11395 14704 11631 14940
rect 11716 14704 11952 14940
rect 12037 14704 12273 14940
rect 12358 14704 12594 14940
rect 12679 14704 12915 14940
rect 13000 14718 13236 14940
rect 13321 14718 13557 14940
rect 13642 14718 13878 14940
rect 13963 14718 14199 14940
rect 13000 14704 13236 14718
rect 13321 14704 13557 14718
rect 13642 14704 13878 14718
rect 13963 14704 14022 14718
rect 14022 14704 14199 14718
rect 14284 14704 14520 14940
rect 14605 14704 14841 14940
rect 9469 14368 9705 14604
rect 9790 14368 10026 14604
rect 10111 14368 10347 14604
rect 10432 14368 10668 14604
rect 10753 14368 10989 14604
rect 11074 14368 11310 14604
rect 11395 14368 11631 14604
rect 11716 14368 11952 14604
rect 12037 14368 12273 14604
rect 12358 14368 12594 14604
rect 12679 14368 12915 14604
rect 13000 14368 13236 14604
rect 13321 14368 13557 14604
rect 13642 14368 13878 14604
rect 13963 14368 14022 14604
rect 14022 14368 14199 14604
rect 14284 14368 14520 14604
rect 14605 14368 14841 14604
rect 9469 14032 9705 14268
rect 9790 14032 10026 14268
rect 10111 14032 10347 14268
rect 10432 14032 10668 14268
rect 10753 14032 10989 14268
rect 11074 14032 11310 14268
rect 11395 14032 11631 14268
rect 11716 14032 11952 14268
rect 12037 14032 12273 14268
rect 12358 14032 12594 14268
rect 12679 14032 12915 14268
rect 13000 14032 13236 14268
rect 13321 14032 13557 14268
rect 13642 14032 13878 14268
rect 13963 14032 14199 14268
rect 14284 14032 14520 14268
rect 14605 14032 14841 14268
<< metal5 >>
rect 0 39965 15000 40000
rect 0 39729 241 39965
rect 477 39729 568 39965
rect 804 39729 895 39965
rect 1131 39729 1222 39965
rect 1458 39729 1549 39965
rect 1785 39729 1876 39965
rect 2112 39729 2203 39965
rect 2439 39729 2530 39965
rect 2766 39729 2857 39965
rect 3093 39729 3184 39965
rect 3420 39729 3511 39965
rect 3747 39729 3838 39965
rect 4074 39729 4165 39965
rect 4401 39729 4492 39965
rect 4728 39729 4819 39965
rect 5055 39729 5146 39965
rect 5382 39729 5473 39965
rect 5709 39729 5800 39965
rect 6036 39729 6127 39965
rect 6363 39729 6454 39965
rect 6690 39729 6781 39965
rect 7017 39729 7108 39965
rect 7344 39729 7435 39965
rect 7671 39729 7762 39965
rect 7998 39729 8089 39965
rect 8325 39729 8415 39965
rect 8651 39729 8741 39965
rect 8977 39729 9067 39965
rect 9303 39729 9393 39965
rect 9629 39729 9719 39965
rect 9955 39729 10045 39965
rect 10281 39729 10371 39965
rect 10607 39729 10697 39965
rect 10933 39729 11023 39965
rect 11259 39729 11349 39965
rect 11585 39729 11675 39965
rect 11911 39729 12001 39965
rect 12237 39729 12327 39965
rect 12563 39729 12653 39965
rect 12889 39729 12979 39965
rect 13215 39729 13305 39965
rect 13541 39729 13631 39965
rect 13867 39729 13957 39965
rect 14193 39729 14283 39965
rect 14519 39729 14609 39965
rect 14845 39729 15000 39965
rect 0 39641 15000 39729
rect 0 39405 241 39641
rect 477 39405 568 39641
rect 804 39405 895 39641
rect 1131 39405 1222 39641
rect 1458 39405 1549 39641
rect 1785 39405 1876 39641
rect 2112 39405 2203 39641
rect 2439 39405 2530 39641
rect 2766 39405 2857 39641
rect 3093 39405 3184 39641
rect 3420 39405 3511 39641
rect 3747 39405 3838 39641
rect 4074 39405 4165 39641
rect 4401 39405 4492 39641
rect 4728 39405 4819 39641
rect 5055 39405 5146 39641
rect 5382 39405 5473 39641
rect 5709 39405 5800 39641
rect 6036 39405 6127 39641
rect 6363 39405 6454 39641
rect 6690 39405 6781 39641
rect 7017 39405 7108 39641
rect 7344 39405 7435 39641
rect 7671 39405 7762 39641
rect 7998 39405 8089 39641
rect 8325 39405 8415 39641
rect 8651 39405 8741 39641
rect 8977 39405 9067 39641
rect 9303 39405 9393 39641
rect 9629 39405 9719 39641
rect 9955 39405 10045 39641
rect 10281 39405 10371 39641
rect 10607 39405 10697 39641
rect 10933 39405 11023 39641
rect 11259 39405 11349 39641
rect 11585 39405 11675 39641
rect 11911 39405 12001 39641
rect 12237 39405 12327 39641
rect 12563 39405 12653 39641
rect 12889 39405 12979 39641
rect 13215 39405 13305 39641
rect 13541 39405 13631 39641
rect 13867 39405 13957 39641
rect 14193 39405 14283 39641
rect 14519 39405 14609 39641
rect 14845 39405 15000 39641
rect 0 39317 15000 39405
rect 0 39081 241 39317
rect 477 39081 568 39317
rect 804 39081 895 39317
rect 1131 39081 1222 39317
rect 1458 39081 1549 39317
rect 1785 39081 1876 39317
rect 2112 39081 2203 39317
rect 2439 39081 2530 39317
rect 2766 39081 2857 39317
rect 3093 39081 3184 39317
rect 3420 39081 3511 39317
rect 3747 39081 3838 39317
rect 4074 39081 4165 39317
rect 4401 39081 4492 39317
rect 4728 39081 4819 39317
rect 5055 39081 5146 39317
rect 5382 39081 5473 39317
rect 5709 39081 5800 39317
rect 6036 39081 6127 39317
rect 6363 39081 6454 39317
rect 6690 39081 6781 39317
rect 7017 39081 7108 39317
rect 7344 39081 7435 39317
rect 7671 39081 7762 39317
rect 7998 39081 8089 39317
rect 8325 39081 8415 39317
rect 8651 39081 8741 39317
rect 8977 39081 9067 39317
rect 9303 39081 9393 39317
rect 9629 39081 9719 39317
rect 9955 39081 10045 39317
rect 10281 39081 10371 39317
rect 10607 39081 10697 39317
rect 10933 39081 11023 39317
rect 11259 39081 11349 39317
rect 11585 39081 11675 39317
rect 11911 39081 12001 39317
rect 12237 39081 12327 39317
rect 12563 39081 12653 39317
rect 12889 39081 12979 39317
rect 13215 39081 13305 39317
rect 13541 39081 13631 39317
rect 13867 39081 13957 39317
rect 14193 39081 14283 39317
rect 14519 39081 14609 39317
rect 14845 39081 15000 39317
rect 0 38993 15000 39081
rect 0 38757 241 38993
rect 477 38757 568 38993
rect 804 38757 895 38993
rect 1131 38757 1222 38993
rect 1458 38757 1549 38993
rect 1785 38757 1876 38993
rect 2112 38757 2203 38993
rect 2439 38757 2530 38993
rect 2766 38757 2857 38993
rect 3093 38757 3184 38993
rect 3420 38757 3511 38993
rect 3747 38757 3838 38993
rect 4074 38757 4165 38993
rect 4401 38757 4492 38993
rect 4728 38757 4819 38993
rect 5055 38757 5146 38993
rect 5382 38757 5473 38993
rect 5709 38757 5800 38993
rect 6036 38757 6127 38993
rect 6363 38757 6454 38993
rect 6690 38757 6781 38993
rect 7017 38757 7108 38993
rect 7344 38757 7435 38993
rect 7671 38757 7762 38993
rect 7998 38757 8089 38993
rect 8325 38757 8415 38993
rect 8651 38757 8741 38993
rect 8977 38757 9067 38993
rect 9303 38757 9393 38993
rect 9629 38757 9719 38993
rect 9955 38757 10045 38993
rect 10281 38757 10371 38993
rect 10607 38757 10697 38993
rect 10933 38757 11023 38993
rect 11259 38757 11349 38993
rect 11585 38757 11675 38993
rect 11911 38757 12001 38993
rect 12237 38757 12327 38993
rect 12563 38757 12653 38993
rect 12889 38757 12979 38993
rect 13215 38757 13305 38993
rect 13541 38757 13631 38993
rect 13867 38757 13957 38993
rect 14193 38757 14283 38993
rect 14519 38757 14609 38993
rect 14845 38757 15000 38993
rect 0 38669 15000 38757
rect 0 38433 241 38669
rect 477 38433 568 38669
rect 804 38433 895 38669
rect 1131 38433 1222 38669
rect 1458 38433 1549 38669
rect 1785 38433 1876 38669
rect 2112 38433 2203 38669
rect 2439 38433 2530 38669
rect 2766 38433 2857 38669
rect 3093 38433 3184 38669
rect 3420 38433 3511 38669
rect 3747 38433 3838 38669
rect 4074 38433 4165 38669
rect 4401 38433 4492 38669
rect 4728 38433 4819 38669
rect 5055 38433 5146 38669
rect 5382 38433 5473 38669
rect 5709 38433 5800 38669
rect 6036 38433 6127 38669
rect 6363 38433 6454 38669
rect 6690 38433 6781 38669
rect 7017 38433 7108 38669
rect 7344 38433 7435 38669
rect 7671 38433 7762 38669
rect 7998 38433 8089 38669
rect 8325 38433 8415 38669
rect 8651 38433 8741 38669
rect 8977 38433 9067 38669
rect 9303 38433 9393 38669
rect 9629 38433 9719 38669
rect 9955 38433 10045 38669
rect 10281 38433 10371 38669
rect 10607 38433 10697 38669
rect 10933 38433 11023 38669
rect 11259 38433 11349 38669
rect 11585 38433 11675 38669
rect 11911 38433 12001 38669
rect 12237 38433 12327 38669
rect 12563 38433 12653 38669
rect 12889 38433 12979 38669
rect 13215 38433 13305 38669
rect 13541 38433 13631 38669
rect 13867 38433 13957 38669
rect 14193 38433 14283 38669
rect 14519 38433 14609 38669
rect 14845 38433 15000 38669
rect 0 38345 15000 38433
rect 0 38109 241 38345
rect 477 38109 568 38345
rect 804 38109 895 38345
rect 1131 38109 1222 38345
rect 1458 38109 1549 38345
rect 1785 38109 1876 38345
rect 2112 38109 2203 38345
rect 2439 38109 2530 38345
rect 2766 38109 2857 38345
rect 3093 38109 3184 38345
rect 3420 38109 3511 38345
rect 3747 38109 3838 38345
rect 4074 38109 4165 38345
rect 4401 38109 4492 38345
rect 4728 38109 4819 38345
rect 5055 38109 5146 38345
rect 5382 38109 5473 38345
rect 5709 38109 5800 38345
rect 6036 38109 6127 38345
rect 6363 38109 6454 38345
rect 6690 38109 6781 38345
rect 7017 38109 7108 38345
rect 7344 38109 7435 38345
rect 7671 38109 7762 38345
rect 7998 38109 8089 38345
rect 8325 38109 8415 38345
rect 8651 38109 8741 38345
rect 8977 38109 9067 38345
rect 9303 38109 9393 38345
rect 9629 38109 9719 38345
rect 9955 38109 10045 38345
rect 10281 38109 10371 38345
rect 10607 38109 10697 38345
rect 10933 38109 11023 38345
rect 11259 38109 11349 38345
rect 11585 38109 11675 38345
rect 11911 38109 12001 38345
rect 12237 38109 12327 38345
rect 12563 38109 12653 38345
rect 12889 38109 12979 38345
rect 13215 38109 13305 38345
rect 13541 38109 13631 38345
rect 13867 38109 13957 38345
rect 14193 38109 14283 38345
rect 14519 38109 14609 38345
rect 14845 38109 15000 38345
rect 0 38021 15000 38109
rect 0 37785 241 38021
rect 477 37785 568 38021
rect 804 37785 895 38021
rect 1131 37785 1222 38021
rect 1458 37785 1549 38021
rect 1785 37785 1876 38021
rect 2112 37785 2203 38021
rect 2439 37785 2530 38021
rect 2766 37785 2857 38021
rect 3093 37785 3184 38021
rect 3420 37785 3511 38021
rect 3747 37785 3838 38021
rect 4074 37785 4165 38021
rect 4401 37785 4492 38021
rect 4728 37785 4819 38021
rect 5055 37785 5146 38021
rect 5382 37785 5473 38021
rect 5709 37785 5800 38021
rect 6036 37785 6127 38021
rect 6363 37785 6454 38021
rect 6690 37785 6781 38021
rect 7017 37785 7108 38021
rect 7344 37785 7435 38021
rect 7671 37785 7762 38021
rect 7998 37785 8089 38021
rect 8325 37785 8415 38021
rect 8651 37785 8741 38021
rect 8977 37785 9067 38021
rect 9303 37785 9393 38021
rect 9629 37785 9719 38021
rect 9955 37785 10045 38021
rect 10281 37785 10371 38021
rect 10607 37785 10697 38021
rect 10933 37785 11023 38021
rect 11259 37785 11349 38021
rect 11585 37785 11675 38021
rect 11911 37785 12001 38021
rect 12237 37785 12327 38021
rect 12563 37785 12653 38021
rect 12889 37785 12979 38021
rect 13215 37785 13305 38021
rect 13541 37785 13631 38021
rect 13867 37785 13957 38021
rect 14193 37785 14283 38021
rect 14519 37785 14609 38021
rect 14845 37785 15000 38021
rect 0 37697 15000 37785
rect 0 37461 241 37697
rect 477 37461 568 37697
rect 804 37461 895 37697
rect 1131 37461 1222 37697
rect 1458 37461 1549 37697
rect 1785 37461 1876 37697
rect 2112 37461 2203 37697
rect 2439 37461 2530 37697
rect 2766 37461 2857 37697
rect 3093 37461 3184 37697
rect 3420 37461 3511 37697
rect 3747 37461 3838 37697
rect 4074 37461 4165 37697
rect 4401 37461 4492 37697
rect 4728 37461 4819 37697
rect 5055 37461 5146 37697
rect 5382 37461 5473 37697
rect 5709 37461 5800 37697
rect 6036 37461 6127 37697
rect 6363 37461 6454 37697
rect 6690 37461 6781 37697
rect 7017 37461 7108 37697
rect 7344 37461 7435 37697
rect 7671 37461 7762 37697
rect 7998 37461 8089 37697
rect 8325 37461 8415 37697
rect 8651 37461 8741 37697
rect 8977 37461 9067 37697
rect 9303 37461 9393 37697
rect 9629 37461 9719 37697
rect 9955 37461 10045 37697
rect 10281 37461 10371 37697
rect 10607 37461 10697 37697
rect 10933 37461 11023 37697
rect 11259 37461 11349 37697
rect 11585 37461 11675 37697
rect 11911 37461 12001 37697
rect 12237 37461 12327 37697
rect 12563 37461 12653 37697
rect 12889 37461 12979 37697
rect 13215 37461 13305 37697
rect 13541 37461 13631 37697
rect 13867 37461 13957 37697
rect 14193 37461 14283 37697
rect 14519 37461 14609 37697
rect 14845 37461 15000 37697
rect 0 37373 15000 37461
rect 0 37137 241 37373
rect 477 37137 568 37373
rect 804 37137 895 37373
rect 1131 37137 1222 37373
rect 1458 37137 1549 37373
rect 1785 37137 1876 37373
rect 2112 37137 2203 37373
rect 2439 37137 2530 37373
rect 2766 37137 2857 37373
rect 3093 37137 3184 37373
rect 3420 37137 3511 37373
rect 3747 37137 3838 37373
rect 4074 37137 4165 37373
rect 4401 37137 4492 37373
rect 4728 37137 4819 37373
rect 5055 37137 5146 37373
rect 5382 37137 5473 37373
rect 5709 37137 5800 37373
rect 6036 37137 6127 37373
rect 6363 37137 6454 37373
rect 6690 37137 6781 37373
rect 7017 37137 7108 37373
rect 7344 37137 7435 37373
rect 7671 37137 7762 37373
rect 7998 37137 8089 37373
rect 8325 37137 8415 37373
rect 8651 37137 8741 37373
rect 8977 37137 9067 37373
rect 9303 37137 9393 37373
rect 9629 37137 9719 37373
rect 9955 37137 10045 37373
rect 10281 37137 10371 37373
rect 10607 37137 10697 37373
rect 10933 37137 11023 37373
rect 11259 37137 11349 37373
rect 11585 37137 11675 37373
rect 11911 37137 12001 37373
rect 12237 37137 12327 37373
rect 12563 37137 12653 37373
rect 12889 37137 12979 37373
rect 13215 37137 13305 37373
rect 13541 37137 13631 37373
rect 13867 37137 13957 37373
rect 14193 37137 14283 37373
rect 14519 37137 14609 37373
rect 14845 37137 15000 37373
rect 0 37049 15000 37137
rect 0 36813 241 37049
rect 477 36813 568 37049
rect 804 36813 895 37049
rect 1131 36813 1222 37049
rect 1458 36813 1549 37049
rect 1785 36813 1876 37049
rect 2112 36813 2203 37049
rect 2439 36813 2530 37049
rect 2766 36813 2857 37049
rect 3093 36813 3184 37049
rect 3420 36813 3511 37049
rect 3747 36813 3838 37049
rect 4074 36813 4165 37049
rect 4401 36813 4492 37049
rect 4728 36813 4819 37049
rect 5055 36813 5146 37049
rect 5382 36813 5473 37049
rect 5709 36813 5800 37049
rect 6036 36813 6127 37049
rect 6363 36813 6454 37049
rect 6690 36813 6781 37049
rect 7017 36813 7108 37049
rect 7344 36813 7435 37049
rect 7671 36813 7762 37049
rect 7998 36813 8089 37049
rect 8325 36813 8415 37049
rect 8651 36813 8741 37049
rect 8977 36813 9067 37049
rect 9303 36813 9393 37049
rect 9629 36813 9719 37049
rect 9955 36813 10045 37049
rect 10281 36813 10371 37049
rect 10607 36813 10697 37049
rect 10933 36813 11023 37049
rect 11259 36813 11349 37049
rect 11585 36813 11675 37049
rect 11911 36813 12001 37049
rect 12237 36813 12327 37049
rect 12563 36813 12653 37049
rect 12889 36813 12979 37049
rect 13215 36813 13305 37049
rect 13541 36813 13631 37049
rect 13867 36813 13957 37049
rect 14193 36813 14283 37049
rect 14519 36813 14609 37049
rect 14845 36813 15000 37049
rect 0 36725 15000 36813
rect 0 36489 241 36725
rect 477 36489 568 36725
rect 804 36489 895 36725
rect 1131 36489 1222 36725
rect 1458 36489 1549 36725
rect 1785 36489 1876 36725
rect 2112 36489 2203 36725
rect 2439 36489 2530 36725
rect 2766 36489 2857 36725
rect 3093 36489 3184 36725
rect 3420 36489 3511 36725
rect 3747 36489 3838 36725
rect 4074 36489 4165 36725
rect 4401 36489 4492 36725
rect 4728 36489 4819 36725
rect 5055 36489 5146 36725
rect 5382 36489 5473 36725
rect 5709 36489 5800 36725
rect 6036 36489 6127 36725
rect 6363 36489 6454 36725
rect 6690 36489 6781 36725
rect 7017 36489 7108 36725
rect 7344 36489 7435 36725
rect 7671 36489 7762 36725
rect 7998 36489 8089 36725
rect 8325 36489 8415 36725
rect 8651 36489 8741 36725
rect 8977 36489 9067 36725
rect 9303 36489 9393 36725
rect 9629 36489 9719 36725
rect 9955 36489 10045 36725
rect 10281 36489 10371 36725
rect 10607 36489 10697 36725
rect 10933 36489 11023 36725
rect 11259 36489 11349 36725
rect 11585 36489 11675 36725
rect 11911 36489 12001 36725
rect 12237 36489 12327 36725
rect 12563 36489 12653 36725
rect 12889 36489 12979 36725
rect 13215 36489 13305 36725
rect 13541 36489 13631 36725
rect 13867 36489 13957 36725
rect 14193 36489 14283 36725
rect 14519 36489 14609 36725
rect 14845 36489 15000 36725
rect 0 36401 15000 36489
rect 0 36165 241 36401
rect 477 36165 568 36401
rect 804 36165 895 36401
rect 1131 36165 1222 36401
rect 1458 36165 1549 36401
rect 1785 36165 1876 36401
rect 2112 36165 2203 36401
rect 2439 36165 2530 36401
rect 2766 36165 2857 36401
rect 3093 36165 3184 36401
rect 3420 36165 3511 36401
rect 3747 36165 3838 36401
rect 4074 36165 4165 36401
rect 4401 36165 4492 36401
rect 4728 36165 4819 36401
rect 5055 36165 5146 36401
rect 5382 36165 5473 36401
rect 5709 36165 5800 36401
rect 6036 36165 6127 36401
rect 6363 36165 6454 36401
rect 6690 36165 6781 36401
rect 7017 36165 7108 36401
rect 7344 36165 7435 36401
rect 7671 36165 7762 36401
rect 7998 36165 8089 36401
rect 8325 36165 8415 36401
rect 8651 36165 8741 36401
rect 8977 36165 9067 36401
rect 9303 36165 9393 36401
rect 9629 36165 9719 36401
rect 9955 36165 10045 36401
rect 10281 36165 10371 36401
rect 10607 36165 10697 36401
rect 10933 36165 11023 36401
rect 11259 36165 11349 36401
rect 11585 36165 11675 36401
rect 11911 36165 12001 36401
rect 12237 36165 12327 36401
rect 12563 36165 12653 36401
rect 12889 36165 12979 36401
rect 13215 36165 13305 36401
rect 13541 36165 13631 36401
rect 13867 36165 13957 36401
rect 14193 36165 14283 36401
rect 14519 36165 14609 36401
rect 14845 36165 15000 36401
rect 0 36077 15000 36165
rect 0 35841 241 36077
rect 477 35841 568 36077
rect 804 35841 895 36077
rect 1131 35841 1222 36077
rect 1458 35841 1549 36077
rect 1785 35841 1876 36077
rect 2112 35841 2203 36077
rect 2439 35841 2530 36077
rect 2766 35841 2857 36077
rect 3093 35841 3184 36077
rect 3420 35841 3511 36077
rect 3747 35841 3838 36077
rect 4074 35841 4165 36077
rect 4401 35841 4492 36077
rect 4728 35841 4819 36077
rect 5055 35841 5146 36077
rect 5382 35841 5473 36077
rect 5709 35841 5800 36077
rect 6036 35841 6127 36077
rect 6363 35841 6454 36077
rect 6690 35841 6781 36077
rect 7017 35841 7108 36077
rect 7344 35841 7435 36077
rect 7671 35841 7762 36077
rect 7998 35841 8089 36077
rect 8325 35841 8415 36077
rect 8651 35841 8741 36077
rect 8977 35841 9067 36077
rect 9303 35841 9393 36077
rect 9629 35841 9719 36077
rect 9955 35841 10045 36077
rect 10281 35841 10371 36077
rect 10607 35841 10697 36077
rect 10933 35841 11023 36077
rect 11259 35841 11349 36077
rect 11585 35841 11675 36077
rect 11911 35841 12001 36077
rect 12237 35841 12327 36077
rect 12563 35841 12653 36077
rect 12889 35841 12979 36077
rect 13215 35841 13305 36077
rect 13541 35841 13631 36077
rect 13867 35841 13957 36077
rect 14193 35841 14283 36077
rect 14519 35841 14609 36077
rect 14845 35841 15000 36077
rect 0 35753 15000 35841
rect 0 35517 241 35753
rect 477 35517 568 35753
rect 804 35517 895 35753
rect 1131 35517 1222 35753
rect 1458 35517 1549 35753
rect 1785 35517 1876 35753
rect 2112 35517 2203 35753
rect 2439 35517 2530 35753
rect 2766 35517 2857 35753
rect 3093 35517 3184 35753
rect 3420 35517 3511 35753
rect 3747 35517 3838 35753
rect 4074 35517 4165 35753
rect 4401 35517 4492 35753
rect 4728 35517 4819 35753
rect 5055 35517 5146 35753
rect 5382 35517 5473 35753
rect 5709 35517 5800 35753
rect 6036 35517 6127 35753
rect 6363 35517 6454 35753
rect 6690 35517 6781 35753
rect 7017 35517 7108 35753
rect 7344 35517 7435 35753
rect 7671 35517 7762 35753
rect 7998 35517 8089 35753
rect 8325 35517 8415 35753
rect 8651 35517 8741 35753
rect 8977 35517 9067 35753
rect 9303 35517 9393 35753
rect 9629 35517 9719 35753
rect 9955 35517 10045 35753
rect 10281 35517 10371 35753
rect 10607 35517 10697 35753
rect 10933 35517 11023 35753
rect 11259 35517 11349 35753
rect 11585 35517 11675 35753
rect 11911 35517 12001 35753
rect 12237 35517 12327 35753
rect 12563 35517 12653 35753
rect 12889 35517 12979 35753
rect 13215 35517 13305 35753
rect 13541 35517 13631 35753
rect 13867 35517 13957 35753
rect 14193 35517 14283 35753
rect 14519 35517 14609 35753
rect 14845 35517 15000 35753
rect 0 35429 15000 35517
rect 0 35193 241 35429
rect 477 35193 568 35429
rect 804 35193 895 35429
rect 1131 35193 1222 35429
rect 1458 35193 1549 35429
rect 1785 35193 1876 35429
rect 2112 35193 2203 35429
rect 2439 35193 2530 35429
rect 2766 35193 2857 35429
rect 3093 35193 3184 35429
rect 3420 35193 3511 35429
rect 3747 35193 3838 35429
rect 4074 35193 4165 35429
rect 4401 35193 4492 35429
rect 4728 35193 4819 35429
rect 5055 35193 5146 35429
rect 5382 35193 5473 35429
rect 5709 35193 5800 35429
rect 6036 35193 6127 35429
rect 6363 35193 6454 35429
rect 6690 35193 6781 35429
rect 7017 35193 7108 35429
rect 7344 35193 7435 35429
rect 7671 35193 7762 35429
rect 7998 35193 8089 35429
rect 8325 35193 8415 35429
rect 8651 35193 8741 35429
rect 8977 35193 9067 35429
rect 9303 35193 9393 35429
rect 9629 35193 9719 35429
rect 9955 35193 10045 35429
rect 10281 35193 10371 35429
rect 10607 35193 10697 35429
rect 10933 35193 11023 35429
rect 11259 35193 11349 35429
rect 11585 35193 11675 35429
rect 11911 35193 12001 35429
rect 12237 35193 12327 35429
rect 12563 35193 12653 35429
rect 12889 35193 12979 35429
rect 13215 35193 13305 35429
rect 13541 35193 13631 35429
rect 13867 35193 13957 35429
rect 14193 35193 14283 35429
rect 14519 35193 14609 35429
rect 14845 35193 15000 35429
rect 0 35157 15000 35193
tri 1933 34288 2265 34620 se
rect 2265 34596 12733 34620
tri 12733 34596 12757 34620 sw
rect 2265 34360 2268 34596
rect 2504 34360 2588 34596
rect 2824 34360 2908 34596
rect 3144 34360 3228 34596
rect 3464 34360 3548 34596
rect 3784 34360 3868 34596
rect 4104 34360 4188 34596
rect 4424 34360 4508 34596
rect 4744 34360 4828 34596
rect 5064 34360 5148 34596
rect 5384 34360 5468 34596
rect 5704 34360 5788 34596
rect 6024 34360 6108 34596
rect 6344 34360 6428 34596
rect 6664 34360 6748 34596
rect 6984 34360 7068 34596
rect 7304 34360 7388 34596
rect 7624 34360 7708 34596
rect 7944 34360 8028 34596
rect 8264 34360 8348 34596
rect 8584 34360 8668 34596
rect 8904 34360 8988 34596
rect 9224 34360 9308 34596
rect 9544 34360 9628 34596
rect 9864 34360 9948 34596
rect 10184 34360 10268 34596
rect 10504 34360 10588 34596
rect 10824 34360 10908 34596
rect 11144 34360 11228 34596
rect 11464 34360 11548 34596
rect 11784 34360 11868 34596
rect 12104 34360 12188 34596
rect 12424 34360 12508 34596
rect 12744 34360 12757 34596
rect 2265 34288 12757 34360
tri 1730 34085 1933 34288 se
rect 1933 34085 1946 34288
tri 1613 33968 1730 34085 se
rect 1730 34052 1946 34085
rect 2182 34234 12757 34288
tri 12757 34234 13119 34596 sw
rect 2182 34232 12870 34234
rect 2182 34212 2404 34232
tri 2404 34212 2424 34232 nw
tri 12577 34212 12597 34232 ne
rect 12597 34212 12870 34232
rect 2182 34197 2389 34212
tri 2389 34197 2404 34212 nw
tri 2417 34197 2432 34212 se
rect 2432 34197 12569 34212
rect 2182 34169 2361 34197
tri 2361 34169 2389 34197 nw
tri 2389 34169 2417 34197 se
rect 2417 34184 12569 34197
tri 12569 34184 12597 34212 sw
tri 12597 34184 12625 34212 ne
rect 12625 34184 12870 34212
rect 2417 34169 12597 34184
rect 2182 34141 2333 34169
tri 2333 34141 2361 34169 nw
tri 2361 34141 2389 34169 se
rect 2389 34156 12597 34169
tri 12597 34156 12625 34184 sw
tri 12625 34156 12653 34184 ne
rect 12653 34156 12870 34184
rect 2389 34141 12625 34156
rect 2182 34113 2305 34141
tri 2305 34113 2333 34141 nw
tri 2333 34113 2361 34141 se
rect 2361 34128 12625 34141
tri 12625 34128 12653 34156 sw
tri 12653 34128 12681 34156 ne
rect 12681 34128 12870 34156
rect 2361 34113 12653 34128
rect 2182 34085 2277 34113
tri 2277 34085 2305 34113 nw
tri 2305 34085 2333 34113 se
rect 2333 34100 12653 34113
tri 12653 34100 12681 34128 sw
tri 12681 34100 12709 34128 ne
rect 12709 34100 12870 34128
rect 2333 34085 12681 34100
rect 2182 34057 2249 34085
tri 2249 34057 2277 34085 nw
tri 2277 34057 2305 34085 se
rect 2305 34072 12681 34085
tri 12681 34072 12709 34100 sw
tri 12709 34072 12737 34100 ne
rect 12737 34072 12870 34100
rect 2305 34057 12709 34072
rect 2182 34052 2221 34057
rect 1730 34029 2221 34052
tri 2221 34029 2249 34057 nw
tri 2249 34029 2277 34057 se
rect 2277 34044 12709 34057
tri 12709 34044 12737 34072 sw
tri 12737 34044 12765 34072 ne
rect 12765 34044 12870 34072
rect 2277 34029 12737 34044
rect 1730 34001 2193 34029
tri 2193 34001 2221 34029 nw
tri 2221 34001 2249 34029 se
rect 2249 34016 12737 34029
tri 12737 34016 12765 34044 sw
tri 12765 34016 12793 34044 ne
rect 12793 34016 12870 34044
rect 2249 34001 12765 34016
rect 1730 33973 2165 34001
tri 2165 33973 2193 34001 nw
tri 2193 33973 2221 34001 se
rect 2221 33988 12765 34001
tri 12765 33988 12793 34016 sw
tri 12793 33988 12821 34016 ne
rect 12821 33998 12870 34016
rect 13106 33998 13119 34234
rect 12821 33988 13119 33998
rect 2221 33973 12793 33988
rect 1730 33968 2137 33973
tri 1293 33648 1613 33968 se
rect 1613 33732 1626 33968
rect 1862 33945 2137 33968
tri 2137 33945 2165 33973 nw
tri 2165 33945 2193 33973 se
rect 2193 33960 12793 33973
tri 12793 33960 12821 33988 sw
tri 12821 33960 12849 33988 ne
rect 12849 33960 13119 33988
rect 2193 33945 12821 33960
rect 1862 33917 2109 33945
tri 2109 33917 2137 33945 nw
tri 2137 33917 2165 33945 se
rect 2165 33932 12821 33945
tri 12821 33932 12849 33960 sw
tri 12849 33932 12877 33960 ne
rect 12877 33932 13119 33960
rect 2165 33917 12849 33932
rect 1862 33889 2081 33917
tri 2081 33889 2109 33917 nw
tri 2109 33889 2137 33917 se
rect 2137 33904 12849 33917
tri 12849 33904 12877 33932 sw
tri 12877 33904 12905 33932 ne
rect 12905 33914 13119 33932
tri 13119 33914 13439 34234 sw
rect 12905 33904 13190 33914
rect 2137 33889 12877 33904
rect 1862 33861 2053 33889
tri 2053 33861 2081 33889 nw
tri 2081 33861 2109 33889 se
rect 2109 33876 12877 33889
tri 12877 33876 12905 33904 sw
tri 12905 33876 12933 33904 ne
rect 12933 33876 13190 33904
rect 2109 33861 12905 33876
rect 1862 33833 2025 33861
tri 2025 33833 2053 33861 nw
tri 2053 33833 2081 33861 se
rect 2081 33848 12905 33861
tri 12905 33848 12933 33876 sw
tri 12933 33848 12961 33876 ne
rect 12961 33848 13190 33876
rect 2081 33833 12933 33848
rect 1862 33805 1997 33833
tri 1997 33805 2025 33833 nw
tri 2025 33805 2053 33833 se
rect 2053 33820 12933 33833
tri 12933 33820 12961 33848 sw
tri 12961 33820 12989 33848 ne
rect 12989 33820 13190 33848
rect 2053 33805 12961 33820
rect 1862 33777 1969 33805
tri 1969 33777 1997 33805 nw
tri 1997 33777 2025 33805 se
rect 2025 33792 12961 33805
tri 12961 33792 12989 33820 sw
tri 12989 33792 13017 33820 ne
rect 13017 33792 13190 33820
rect 2025 33777 12989 33792
rect 1862 33749 1941 33777
tri 1941 33749 1969 33777 nw
tri 1969 33749 1997 33777 se
rect 1997 33764 12989 33777
tri 12989 33764 13017 33792 sw
tri 13017 33764 13045 33792 ne
rect 13045 33764 13190 33792
rect 1997 33749 13017 33764
rect 1862 33732 1913 33749
rect 1613 33721 1913 33732
tri 1913 33721 1941 33749 nw
tri 1941 33721 1969 33749 se
rect 1969 33736 13017 33749
tri 13017 33736 13045 33764 sw
tri 13045 33736 13073 33764 ne
rect 13073 33736 13190 33764
rect 1969 33721 13045 33736
rect 1613 33693 1885 33721
tri 1885 33693 1913 33721 nw
tri 1913 33693 1941 33721 se
rect 1941 33708 13045 33721
tri 13045 33708 13073 33736 sw
tri 13073 33708 13101 33736 ne
rect 13101 33708 13190 33736
rect 1941 33693 13073 33708
rect 1613 33665 1857 33693
tri 1857 33665 1885 33693 nw
tri 1885 33665 1913 33693 se
rect 1913 33680 13073 33693
tri 13073 33680 13101 33708 sw
tri 13101 33680 13129 33708 ne
rect 13129 33680 13190 33708
rect 1913 33665 13101 33680
rect 1613 33648 1829 33665
tri 1198 33553 1293 33648 se
rect 1293 33553 1306 33648
tri 970 33325 1198 33553 se
rect 1198 33412 1306 33553
rect 1542 33637 1829 33648
tri 1829 33637 1857 33665 nw
tri 1857 33637 1885 33665 se
rect 1885 33652 13101 33665
tri 13101 33652 13129 33680 sw
tri 13129 33652 13157 33680 ne
rect 13157 33678 13190 33680
rect 13426 33678 13439 33914
rect 13157 33652 13439 33678
rect 1885 33637 13129 33652
rect 1542 33609 1801 33637
tri 1801 33609 1829 33637 nw
tri 1829 33609 1857 33637 se
rect 1857 33624 13129 33637
tri 13129 33624 13157 33652 sw
tri 13157 33624 13185 33652 ne
rect 13185 33624 13439 33652
rect 1857 33609 13157 33624
rect 1542 33581 1773 33609
tri 1773 33581 1801 33609 nw
tri 1801 33581 1829 33609 se
rect 1829 33596 13157 33609
tri 13157 33596 13185 33624 sw
tri 13185 33596 13213 33624 ne
rect 13213 33596 13439 33624
rect 1829 33581 13185 33596
rect 1542 33553 1745 33581
tri 1745 33553 1773 33581 nw
tri 1773 33553 1801 33581 se
rect 1801 33568 13185 33581
tri 13185 33568 13213 33596 sw
tri 13213 33568 13241 33596 ne
rect 13241 33594 13439 33596
tri 13439 33594 13759 33914 sw
rect 13241 33568 13510 33594
rect 1801 33553 13213 33568
rect 1542 33525 1717 33553
tri 1717 33525 1745 33553 nw
tri 1745 33525 1773 33553 se
rect 1773 33540 13213 33553
tri 13213 33540 13241 33568 sw
tri 13241 33540 13269 33568 ne
rect 13269 33540 13510 33568
rect 1773 33525 13241 33540
rect 1542 33497 1689 33525
tri 1689 33497 1717 33525 nw
tri 1717 33497 1745 33525 se
rect 1745 33512 13241 33525
tri 13241 33512 13269 33540 sw
tri 13269 33512 13297 33540 ne
rect 13297 33512 13510 33540
rect 1745 33497 13269 33512
rect 1542 33469 1661 33497
tri 1661 33469 1689 33497 nw
tri 1689 33469 1717 33497 se
rect 1717 33484 13269 33497
tri 13269 33484 13297 33512 sw
tri 13297 33484 13325 33512 ne
rect 13325 33484 13510 33512
rect 1717 33469 13297 33484
rect 1542 33441 1633 33469
tri 1633 33441 1661 33469 nw
tri 1661 33441 1689 33469 se
rect 1689 33456 13297 33469
tri 13297 33456 13325 33484 sw
tri 13325 33456 13353 33484 ne
rect 13353 33456 13510 33484
rect 1689 33441 13325 33456
rect 1542 33413 1605 33441
tri 1605 33413 1633 33441 nw
tri 1633 33413 1661 33441 se
rect 1661 33428 13325 33441
tri 13325 33428 13353 33456 sw
tri 13353 33428 13381 33456 ne
rect 13381 33428 13510 33456
rect 1661 33413 13353 33428
rect 1542 33412 1577 33413
rect 1198 33385 1577 33412
tri 1577 33385 1605 33413 nw
tri 1605 33385 1633 33413 se
rect 1633 33400 13353 33413
tri 13353 33400 13381 33428 sw
tri 13381 33400 13409 33428 ne
rect 13409 33400 13510 33428
rect 1633 33385 13381 33400
rect 1198 33357 1549 33385
tri 1549 33357 1577 33385 nw
tri 1577 33357 1605 33385 se
rect 1605 33372 13381 33385
tri 13381 33372 13409 33400 sw
tri 13409 33372 13437 33400 ne
rect 13437 33372 13510 33400
rect 1605 33357 13409 33372
rect 1198 33329 1521 33357
tri 1521 33329 1549 33357 nw
tri 1549 33329 1577 33357 se
rect 1577 33344 13409 33357
tri 13409 33344 13437 33372 sw
tri 13437 33344 13465 33372 ne
rect 13465 33358 13510 33372
rect 13746 33358 13759 33594
rect 13465 33344 13759 33358
rect 1577 33329 13437 33344
rect 1198 33325 1493 33329
tri 959 33314 970 33325 se
rect 970 33314 983 33325
rect 959 33089 983 33314
rect 1219 33301 1493 33325
tri 1493 33301 1521 33329 nw
tri 1521 33301 1549 33329 se
rect 1549 33316 13437 33329
tri 13437 33316 13465 33344 sw
tri 13465 33316 13493 33344 ne
rect 13493 33316 13759 33344
rect 1549 33301 13465 33316
rect 1219 33273 1465 33301
tri 1465 33273 1493 33301 nw
tri 1493 33273 1521 33301 se
rect 1521 33288 13465 33301
tri 13465 33288 13493 33316 sw
tri 13493 33288 13521 33316 ne
rect 13521 33314 13759 33316
tri 13759 33314 14039 33594 sw
rect 13521 33288 14039 33314
rect 1521 33273 13493 33288
rect 1219 33245 1437 33273
tri 1437 33245 1465 33273 nw
tri 1465 33245 1493 33273 se
rect 1493 33260 13493 33273
tri 13493 33260 13521 33288 sw
tri 13521 33260 13549 33288 ne
rect 13549 33260 14039 33288
rect 1493 33245 13521 33260
rect 1219 33217 1409 33245
tri 1409 33217 1437 33245 nw
tri 1437 33217 1465 33245 se
rect 1465 33232 13521 33245
tri 13521 33232 13549 33260 sw
tri 13549 33232 13577 33260 ne
rect 13577 33232 14039 33260
rect 1465 33217 13549 33232
rect 1219 33189 1381 33217
tri 1381 33189 1409 33217 nw
tri 1409 33189 1437 33217 se
rect 1437 33204 13549 33217
tri 13549 33204 13577 33232 sw
tri 13577 33204 13605 33232 ne
rect 13605 33231 14039 33232
rect 13605 33204 13779 33231
rect 1437 33189 13577 33204
rect 1219 33161 1353 33189
tri 1353 33161 1381 33189 nw
tri 1381 33161 1409 33189 se
rect 1409 33178 13577 33189
tri 13577 33178 13603 33204 sw
tri 13605 33186 13623 33204 ne
rect 1409 33161 13603 33178
rect 1219 33089 1333 33161
tri 1333 33141 1353 33161 nw
rect 959 33005 1333 33089
rect 959 32769 983 33005
rect 1219 32769 1333 33005
rect 959 32685 1333 32769
rect 959 32449 983 32685
rect 1219 32449 1333 32685
rect 959 32365 1333 32449
rect 959 32129 983 32365
rect 1219 32129 1333 32365
rect 959 32045 1333 32129
rect 959 31809 983 32045
rect 1219 31809 1333 32045
rect 959 31725 1333 31809
rect 959 31489 983 31725
rect 1219 31489 1333 31725
rect 959 31405 1333 31489
rect 959 31169 983 31405
rect 1219 31169 1333 31405
rect 959 31085 1333 31169
rect 959 30849 983 31085
rect 1219 30849 1333 31085
rect 959 30765 1333 30849
rect 959 30529 983 30765
rect 1219 30529 1333 30765
rect 959 30445 1333 30529
rect 959 30209 983 30445
rect 1219 30209 1333 30445
rect 959 30125 1333 30209
rect 959 29889 983 30125
rect 1219 29889 1333 30125
rect 959 29805 1333 29889
rect 959 29569 983 29805
rect 1219 29569 1333 29805
rect 959 29485 1333 29569
rect 959 29249 983 29485
rect 1219 29249 1333 29485
rect 959 29165 1333 29249
rect 959 28929 983 29165
rect 1219 28929 1333 29165
rect 959 28845 1333 28929
rect 959 28609 983 28845
rect 1219 28609 1333 28845
rect 959 28525 1333 28609
rect 959 28289 983 28525
rect 1219 28289 1333 28525
rect 959 28205 1333 28289
rect 959 27969 983 28205
rect 1219 27969 1333 28205
rect 959 27885 1333 27969
rect 959 27649 983 27885
rect 1219 27649 1333 27885
rect 959 27565 1333 27649
rect 959 27329 983 27565
rect 1219 27329 1333 27565
rect 959 27245 1333 27329
rect 959 27009 983 27245
rect 1219 27009 1333 27245
rect 959 26925 1333 27009
rect 959 26689 983 26925
rect 1219 26689 1333 26925
rect 959 26605 1333 26689
rect 959 26369 983 26605
rect 1219 26369 1333 26605
rect 959 26285 1333 26369
rect 959 26049 983 26285
rect 1219 26049 1333 26285
rect 959 25965 1333 26049
rect 959 25729 983 25965
rect 1219 25729 1333 25965
rect 959 25645 1333 25729
rect 959 25409 983 25645
rect 1219 25409 1333 25645
rect 959 25325 1333 25409
rect 959 25089 983 25325
rect 1219 25089 1333 25325
rect 959 25005 1333 25089
rect 959 24769 983 25005
rect 1219 24769 1333 25005
rect 959 24685 1333 24769
rect 959 24449 983 24685
rect 1219 24449 1333 24685
rect 959 24365 1333 24449
rect 959 24129 983 24365
rect 1219 24129 1333 24365
rect 959 24045 1333 24129
rect 959 23809 983 24045
rect 1219 23809 1333 24045
rect 959 23725 1333 23809
rect 959 23489 983 23725
rect 1219 23489 1333 23725
rect 959 23405 1333 23489
rect 959 23169 983 23405
rect 1219 23169 1333 23405
rect 959 23085 1333 23169
rect 959 22849 983 23085
rect 1219 22849 1333 23085
rect 959 22765 1333 22849
rect 959 22529 983 22765
rect 1219 22529 1333 22765
rect 959 22445 1333 22529
rect 959 22209 983 22445
rect 1219 22209 1333 22445
rect 959 22125 1333 22209
rect 959 21889 983 22125
rect 1219 21889 1333 22125
rect 959 21805 1333 21889
rect 959 21569 983 21805
rect 1219 21569 1333 21805
rect 959 21485 1333 21569
rect 959 21249 983 21485
rect 1219 21249 1333 21485
rect 959 21165 1333 21249
rect 959 20929 983 21165
rect 1219 21049 1333 21165
tri 1353 33133 1381 33161 se
rect 1381 33133 13603 33161
rect 1353 21077 13603 33133
tri 1333 21049 1353 21069 sw
tri 1353 21049 1381 21077 ne
rect 1381 21049 13603 21077
rect 1219 21024 1353 21049
tri 1353 21024 1378 21049 sw
tri 1381 21024 1406 21049 ne
rect 1406 21024 13603 21049
rect 1219 20996 1378 21024
tri 1378 20996 1406 21024 sw
tri 1406 20996 1434 21024 ne
rect 1434 21022 13603 21024
rect 1434 20996 13575 21022
rect 1219 20968 1406 20996
tri 1406 20968 1434 20996 sw
tri 1434 20968 1462 20996 ne
rect 1462 20994 13575 20996
tri 13575 20994 13603 21022 nw
rect 13623 32995 13779 33204
rect 14015 32995 14039 33231
rect 13623 32911 14039 32995
rect 13623 32675 13779 32911
rect 14015 32675 14039 32911
rect 13623 32591 14039 32675
rect 13623 32355 13779 32591
rect 14015 32355 14039 32591
rect 13623 32271 14039 32355
rect 13623 32035 13779 32271
rect 14015 32035 14039 32271
rect 13623 31951 14039 32035
rect 13623 31715 13779 31951
rect 14015 31715 14039 31951
rect 13623 31631 14039 31715
rect 13623 31395 13779 31631
rect 14015 31395 14039 31631
rect 13623 31311 14039 31395
rect 13623 31075 13779 31311
rect 14015 31075 14039 31311
rect 13623 30991 14039 31075
rect 13623 30755 13779 30991
rect 14015 30755 14039 30991
rect 13623 30671 14039 30755
rect 13623 30435 13779 30671
rect 14015 30435 14039 30671
rect 13623 30351 14039 30435
rect 13623 30115 13779 30351
rect 14015 30115 14039 30351
rect 13623 30031 14039 30115
rect 13623 29795 13779 30031
rect 14015 29795 14039 30031
rect 13623 29711 14039 29795
rect 13623 29475 13779 29711
rect 14015 29475 14039 29711
rect 13623 29391 14039 29475
rect 13623 29155 13779 29391
rect 14015 29155 14039 29391
rect 13623 29071 14039 29155
rect 13623 28835 13779 29071
rect 14015 28835 14039 29071
rect 13623 28751 14039 28835
rect 13623 28515 13779 28751
rect 14015 28515 14039 28751
rect 13623 28431 14039 28515
rect 13623 28195 13779 28431
rect 14015 28195 14039 28431
rect 13623 28111 14039 28195
rect 13623 27875 13779 28111
rect 14015 27875 14039 28111
rect 13623 27791 14039 27875
rect 13623 27555 13779 27791
rect 14015 27555 14039 27791
rect 13623 27471 14039 27555
rect 13623 27235 13779 27471
rect 14015 27235 14039 27471
rect 13623 27151 14039 27235
rect 13623 26915 13779 27151
rect 14015 26915 14039 27151
rect 13623 26831 14039 26915
rect 13623 26595 13779 26831
rect 14015 26595 14039 26831
rect 13623 26511 14039 26595
rect 13623 26275 13779 26511
rect 14015 26275 14039 26511
rect 13623 26191 14039 26275
rect 13623 25955 13779 26191
rect 14015 25955 14039 26191
rect 13623 25871 14039 25955
rect 13623 25635 13779 25871
rect 14015 25635 14039 25871
rect 13623 25551 14039 25635
rect 13623 25315 13779 25551
rect 14015 25315 14039 25551
rect 13623 25231 14039 25315
rect 13623 24995 13779 25231
rect 14015 24995 14039 25231
rect 13623 24911 14039 24995
rect 13623 24675 13779 24911
rect 14015 24675 14039 24911
rect 13623 24591 14039 24675
rect 13623 24355 13779 24591
rect 14015 24355 14039 24591
rect 13623 24271 14039 24355
rect 13623 24035 13779 24271
rect 14015 24035 14039 24271
rect 13623 23951 14039 24035
rect 13623 23715 13779 23951
rect 14015 23715 14039 23951
rect 13623 23631 14039 23715
rect 13623 23395 13779 23631
rect 14015 23395 14039 23631
rect 13623 23311 14039 23395
rect 13623 23075 13779 23311
rect 14015 23075 14039 23311
rect 13623 22991 14039 23075
rect 13623 22755 13779 22991
rect 14015 22755 14039 22991
rect 13623 22671 14039 22755
rect 13623 22435 13779 22671
rect 14015 22435 14039 22671
rect 13623 22351 14039 22435
rect 13623 22115 13779 22351
rect 14015 22115 14039 22351
rect 13623 22031 14039 22115
rect 13623 21795 13779 22031
rect 14015 21795 14039 22031
rect 13623 21711 14039 21795
rect 13623 21475 13779 21711
rect 14015 21475 14039 21711
rect 13623 21391 14039 21475
rect 13623 21155 13779 21391
rect 14015 21155 14039 21391
rect 13623 21071 14039 21155
tri 13603 20994 13623 21014 se
rect 13623 20994 13779 21071
rect 1462 20968 13547 20994
rect 1219 20940 1434 20968
tri 1434 20940 1462 20968 sw
tri 1462 20940 1490 20968 ne
rect 1490 20966 13547 20968
tri 13547 20966 13575 20994 nw
tri 13575 20966 13603 20994 se
rect 13603 20966 13779 20994
rect 1490 20940 13519 20966
rect 1219 20929 1462 20940
rect 959 20912 1462 20929
tri 1462 20912 1490 20940 sw
tri 1490 20912 1518 20940 ne
rect 1518 20938 13519 20940
tri 13519 20938 13547 20966 nw
tri 13547 20938 13575 20966 se
rect 13575 20938 13779 20966
rect 1518 20912 13491 20938
rect 959 20884 1490 20912
tri 1490 20884 1518 20912 sw
tri 1518 20884 1546 20912 ne
rect 1546 20910 13491 20912
tri 13491 20910 13519 20938 nw
tri 13519 20910 13547 20938 se
rect 13547 20910 13779 20938
rect 1546 20884 13463 20910
rect 959 20856 1518 20884
tri 1518 20856 1546 20884 sw
tri 1546 20856 1574 20884 ne
rect 1574 20882 13463 20884
tri 13463 20882 13491 20910 nw
tri 13491 20882 13519 20910 se
rect 13519 20882 13779 20910
rect 1574 20856 13435 20882
rect 959 20846 1546 20856
tri 959 20566 1239 20846 ne
rect 1239 20828 1546 20846
tri 1546 20828 1574 20856 sw
tri 1574 20828 1602 20856 ne
rect 1602 20854 13435 20856
tri 13435 20854 13463 20882 nw
tri 13463 20854 13491 20882 se
rect 13491 20854 13779 20882
rect 1602 20828 13407 20854
rect 1239 20802 1574 20828
rect 1239 20566 1252 20802
rect 1488 20800 1574 20802
tri 1574 20800 1602 20828 sw
tri 1602 20800 1630 20828 ne
rect 1630 20826 13407 20828
tri 13407 20826 13435 20854 nw
tri 13435 20826 13463 20854 se
rect 13463 20835 13779 20854
rect 14015 20846 14039 21071
rect 14015 20835 14019 20846
rect 13463 20826 14019 20835
tri 14019 20826 14039 20846 nw
rect 1630 20800 13379 20826
rect 1488 20772 1602 20800
tri 1602 20772 1630 20800 sw
tri 1630 20772 1658 20800 ne
rect 1658 20798 13379 20800
tri 13379 20798 13407 20826 nw
tri 13407 20798 13435 20826 se
rect 13435 20798 13705 20826
rect 1658 20772 13351 20798
rect 1488 20744 1630 20772
tri 1630 20744 1658 20772 sw
tri 1658 20744 1686 20772 ne
rect 1686 20770 13351 20772
tri 13351 20770 13379 20798 nw
tri 13379 20770 13407 20798 se
rect 13407 20770 13705 20798
rect 1686 20744 13323 20770
rect 1488 20716 1658 20744
tri 1658 20716 1686 20744 sw
tri 1686 20716 1714 20744 ne
rect 1714 20742 13323 20744
tri 13323 20742 13351 20770 nw
tri 13351 20742 13379 20770 se
rect 13379 20748 13705 20770
rect 13379 20742 13456 20748
rect 1714 20716 13295 20742
rect 1488 20688 1686 20716
tri 1686 20688 1714 20716 sw
tri 1714 20688 1742 20716 ne
rect 1742 20714 13295 20716
tri 13295 20714 13323 20742 nw
tri 13323 20714 13351 20742 se
rect 13351 20714 13456 20742
rect 1742 20688 13267 20714
rect 1488 20660 1714 20688
tri 1714 20660 1742 20688 sw
tri 1742 20660 1770 20688 ne
rect 1770 20686 13267 20688
tri 13267 20686 13295 20714 nw
tri 13295 20686 13323 20714 se
rect 13323 20686 13456 20714
rect 1770 20660 13239 20686
rect 1488 20632 1742 20660
tri 1742 20632 1770 20660 sw
tri 1770 20632 1798 20660 ne
rect 1798 20658 13239 20660
tri 13239 20658 13267 20686 nw
tri 13267 20658 13295 20686 se
rect 13295 20658 13456 20686
rect 1798 20632 13211 20658
rect 1488 20604 1770 20632
tri 1770 20604 1798 20632 sw
tri 1798 20604 1826 20632 ne
rect 1826 20630 13211 20632
tri 13211 20630 13239 20658 nw
tri 13239 20630 13267 20658 se
rect 13267 20630 13456 20658
rect 1826 20604 13183 20630
rect 1488 20576 1798 20604
tri 1798 20576 1826 20604 sw
tri 1826 20576 1854 20604 ne
rect 1854 20602 13183 20604
tri 13183 20602 13211 20630 nw
tri 13211 20602 13239 20630 se
rect 13239 20602 13456 20630
rect 1854 20576 13155 20602
rect 1488 20566 1826 20576
tri 1239 20240 1565 20566 ne
rect 1565 20548 1826 20566
tri 1826 20548 1854 20576 sw
tri 1854 20548 1882 20576 ne
rect 1882 20574 13155 20576
tri 13155 20574 13183 20602 nw
tri 13183 20574 13211 20602 se
rect 13211 20574 13456 20602
rect 1882 20548 13127 20574
rect 1565 20520 1854 20548
tri 1854 20520 1882 20548 sw
tri 1882 20520 1910 20548 ne
rect 1910 20546 13127 20548
tri 13127 20546 13155 20574 nw
tri 13155 20546 13183 20574 se
rect 13183 20546 13456 20574
rect 1910 20520 13099 20546
rect 1565 20492 1882 20520
tri 1882 20492 1910 20520 sw
tri 1910 20492 1938 20520 ne
rect 1938 20518 13099 20520
tri 13099 20518 13127 20546 nw
tri 13127 20518 13155 20546 se
rect 13155 20518 13456 20546
rect 1938 20492 13071 20518
rect 1565 20482 1910 20492
rect 1565 20246 1572 20482
rect 1808 20464 1910 20482
tri 1910 20464 1938 20492 sw
tri 1938 20464 1966 20492 ne
rect 1966 20490 13071 20492
tri 13071 20490 13099 20518 nw
tri 13099 20490 13127 20518 se
rect 13127 20512 13456 20518
rect 13692 20512 13705 20748
tri 13705 20512 14019 20826 nw
rect 13127 20490 13375 20512
rect 1966 20464 13043 20490
rect 1808 20436 1938 20464
tri 1938 20436 1966 20464 sw
tri 1966 20436 1994 20464 ne
rect 1994 20462 13043 20464
tri 13043 20462 13071 20490 nw
tri 13071 20462 13099 20490 se
rect 13099 20462 13375 20490
rect 1994 20436 13015 20462
rect 1808 20408 1966 20436
tri 1966 20408 1994 20436 sw
tri 1994 20408 2022 20436 ne
rect 2022 20434 13015 20436
tri 13015 20434 13043 20462 nw
tri 13043 20434 13071 20462 se
rect 13071 20434 13375 20462
rect 2022 20408 12987 20434
rect 1808 20380 1994 20408
tri 1994 20380 2022 20408 sw
tri 2022 20380 2050 20408 ne
rect 2050 20406 12987 20408
tri 12987 20406 13015 20434 nw
tri 13015 20406 13043 20434 se
rect 13043 20428 13375 20434
rect 13043 20406 13136 20428
rect 2050 20380 12959 20406
rect 1808 20352 2022 20380
tri 2022 20352 2050 20380 sw
tri 2050 20352 2078 20380 ne
rect 2078 20378 12959 20380
tri 12959 20378 12987 20406 nw
tri 12987 20378 13015 20406 se
rect 13015 20378 13136 20406
rect 2078 20352 12931 20378
rect 1808 20324 2050 20352
tri 2050 20324 2078 20352 sw
tri 2078 20324 2106 20352 ne
rect 2106 20350 12931 20352
tri 12931 20350 12959 20378 nw
tri 12959 20350 12987 20378 se
rect 12987 20350 13136 20378
rect 2106 20324 12903 20350
rect 1808 20296 2078 20324
tri 2078 20296 2106 20324 sw
tri 2106 20296 2134 20324 ne
rect 2134 20322 12903 20324
tri 12903 20322 12931 20350 nw
tri 12931 20322 12959 20350 se
rect 12959 20322 13136 20350
rect 2134 20296 12875 20322
rect 1808 20268 2106 20296
tri 2106 20268 2134 20296 sw
tri 2134 20268 2162 20296 ne
rect 2162 20294 12875 20296
tri 12875 20294 12903 20322 nw
tri 12903 20294 12931 20322 se
rect 12931 20294 13136 20322
rect 2162 20268 12847 20294
rect 1808 20246 2134 20268
rect 1565 20240 2134 20246
tri 2134 20240 2162 20268 sw
tri 2162 20240 2190 20268 ne
rect 2190 20266 12847 20268
tri 12847 20266 12875 20294 nw
tri 12875 20266 12903 20294 se
rect 12903 20266 13136 20294
rect 2190 20240 12819 20266
tri 1565 19926 1879 20240 ne
rect 1879 20212 2162 20240
tri 2162 20212 2190 20240 sw
tri 2190 20212 2218 20240 ne
rect 2218 20238 12819 20240
tri 12819 20238 12847 20266 nw
tri 12847 20238 12875 20266 se
rect 12875 20238 13136 20266
rect 2218 20212 12791 20238
rect 1879 20184 2190 20212
tri 2190 20184 2218 20212 sw
tri 2218 20184 2246 20212 ne
rect 2246 20210 12791 20212
tri 12791 20210 12819 20238 nw
tri 12819 20210 12847 20238 se
rect 12847 20210 13136 20238
rect 2246 20184 12763 20210
rect 1879 20162 2218 20184
rect 1879 19926 1892 20162
rect 2128 20156 2218 20162
tri 2218 20156 2246 20184 sw
tri 2246 20156 2274 20184 ne
rect 2274 20182 12763 20184
tri 12763 20182 12791 20210 nw
tri 12791 20182 12819 20210 se
rect 12819 20192 13136 20210
rect 13372 20192 13375 20428
rect 12819 20182 13375 20192
tri 13375 20182 13705 20512 nw
rect 2274 20156 12735 20182
rect 2128 20128 2246 20156
tri 2246 20128 2274 20156 sw
tri 2274 20128 2302 20156 ne
rect 2302 20154 12735 20156
tri 12735 20154 12763 20182 nw
tri 12763 20154 12791 20182 se
rect 12791 20154 13065 20182
rect 2302 20128 12707 20154
rect 2128 20100 2274 20128
tri 2274 20100 2302 20128 sw
tri 2302 20100 2330 20128 ne
rect 2330 20126 12707 20128
tri 12707 20126 12735 20154 nw
tri 12735 20126 12763 20154 se
rect 12763 20126 13065 20154
rect 2330 20100 12679 20126
rect 2128 20072 2302 20100
tri 2302 20072 2330 20100 sw
tri 2330 20072 2358 20100 ne
rect 2358 20098 12679 20100
tri 12679 20098 12707 20126 nw
tri 12707 20098 12735 20126 se
rect 12735 20108 13065 20126
rect 12735 20098 12816 20108
rect 2358 20072 12651 20098
rect 2128 20044 2330 20072
tri 2330 20044 2358 20072 sw
tri 2358 20044 2386 20072 ne
rect 2386 20070 12651 20072
tri 12651 20070 12679 20098 nw
tri 12679 20070 12707 20098 se
rect 12707 20070 12816 20098
rect 2386 20044 12623 20070
rect 2128 20016 2358 20044
tri 2358 20016 2386 20044 sw
tri 2386 20016 2414 20044 ne
rect 2414 20042 12623 20044
tri 12623 20042 12651 20070 nw
tri 12651 20042 12679 20070 se
rect 12679 20042 12816 20070
rect 2414 20016 12595 20042
rect 2128 19988 2386 20016
tri 2386 19988 2414 20016 sw
tri 2414 19988 2442 20016 ne
rect 2442 20014 12595 20016
tri 12595 20014 12623 20042 nw
tri 12623 20014 12651 20042 se
rect 12651 20014 12816 20042
rect 2442 19988 12567 20014
rect 2128 19960 2414 19988
tri 2414 19960 2442 19988 sw
tri 2442 19960 2470 19988 ne
rect 2470 19986 12567 19988
tri 12567 19986 12595 20014 nw
tri 12595 19986 12623 20014 se
rect 12623 19986 12816 20014
rect 2470 19960 12539 19986
rect 2128 19932 2442 19960
tri 2442 19932 2470 19960 sw
tri 2470 19932 2498 19960 ne
rect 2498 19958 12539 19960
tri 12539 19958 12567 19986 nw
tri 12567 19958 12595 19986 se
rect 12595 19958 12816 19986
rect 2498 19932 12511 19958
rect 2128 19926 2470 19932
tri 1879 19564 2241 19926 ne
rect 2241 19904 2470 19926
tri 2470 19904 2498 19932 sw
tri 2498 19904 2526 19932 ne
rect 2526 19930 12511 19932
tri 12511 19930 12539 19958 nw
tri 12539 19930 12567 19958 se
rect 12567 19930 12816 19958
rect 2526 19904 12485 19930
tri 12485 19904 12511 19930 nw
tri 12513 19904 12539 19930 se
rect 12539 19904 12816 19930
rect 2241 19884 2498 19904
tri 2498 19884 2518 19904 sw
tri 12493 19884 12513 19904 se
rect 12513 19884 12816 19904
rect 2241 19872 12816 19884
rect 13052 19872 13065 20108
tri 13065 19872 13375 20182 nw
rect 2241 19800 12733 19872
rect 2241 19564 2254 19800
rect 2490 19564 2574 19800
rect 2810 19564 2894 19800
rect 3130 19564 3214 19800
rect 3450 19564 3534 19800
rect 3770 19564 3854 19800
rect 4090 19564 4174 19800
rect 4410 19564 4494 19800
rect 4730 19564 4814 19800
rect 5050 19564 5134 19800
rect 5370 19564 5454 19800
rect 5690 19564 5774 19800
rect 6010 19564 6094 19800
rect 6330 19564 6414 19800
rect 6650 19564 6734 19800
rect 6970 19564 7054 19800
rect 7290 19564 7374 19800
rect 7610 19564 7694 19800
rect 7930 19564 8014 19800
rect 8250 19564 8334 19800
rect 8570 19564 8654 19800
rect 8890 19564 8974 19800
rect 9210 19564 9294 19800
rect 9530 19564 9614 19800
rect 9850 19564 9934 19800
rect 10170 19564 10254 19800
rect 10490 19564 10574 19800
rect 10810 19564 10894 19800
rect 11130 19564 11214 19800
rect 11450 19564 11534 19800
rect 11770 19564 11854 19800
rect 12090 19564 12174 19800
rect 12410 19564 12494 19800
rect 12730 19564 12733 19800
tri 2241 19540 2265 19564 ne
rect 2265 19540 12733 19564
tri 12733 19540 13065 19872 nw
rect 0 18972 15000 18997
rect 0 18736 143 18972
rect 379 18736 465 18972
rect 701 18736 787 18972
rect 1023 18736 1109 18972
rect 1345 18736 1431 18972
rect 1667 18736 1753 18972
rect 1989 18736 2075 18972
rect 2311 18736 2397 18972
rect 2633 18736 2719 18972
rect 2955 18736 3041 18972
rect 3277 18736 3363 18972
rect 3599 18736 3685 18972
rect 3921 18736 4007 18972
rect 4243 18736 4329 18972
rect 4565 18736 4651 18972
rect 4887 18736 4973 18972
rect 5209 18736 5295 18972
rect 5531 18736 9469 18972
rect 9705 18736 9790 18972
rect 10026 18736 10111 18972
rect 10347 18736 10432 18972
rect 10668 18736 10753 18972
rect 10989 18736 11074 18972
rect 11310 18736 11395 18972
rect 11631 18736 11716 18972
rect 11952 18736 12037 18972
rect 12273 18736 12358 18972
rect 12594 18736 12679 18972
rect 12915 18736 13000 18972
rect 13236 18736 13321 18972
rect 13557 18736 13642 18972
rect 13878 18736 13963 18972
rect 14199 18736 14284 18972
rect 14520 18736 14605 18972
rect 14841 18736 15000 18972
rect 0 18636 15000 18736
rect 0 18400 143 18636
rect 379 18400 465 18636
rect 701 18400 787 18636
rect 1023 18400 1109 18636
rect 1345 18400 1431 18636
rect 1667 18400 1753 18636
rect 1989 18400 2075 18636
rect 2311 18400 2397 18636
rect 2633 18400 2719 18636
rect 2955 18400 3041 18636
rect 3277 18400 3363 18636
rect 3599 18400 3685 18636
rect 3921 18400 4007 18636
rect 4243 18400 4329 18636
rect 4565 18400 4651 18636
rect 4887 18400 4973 18636
rect 5209 18400 5295 18636
rect 5531 18400 9469 18636
rect 9705 18400 9790 18636
rect 10026 18400 10111 18636
rect 10347 18400 10432 18636
rect 10668 18400 10753 18636
rect 10989 18400 11074 18636
rect 11310 18400 11395 18636
rect 11631 18400 11716 18636
rect 11952 18400 12037 18636
rect 12273 18400 12358 18636
rect 12594 18400 12679 18636
rect 12915 18400 13000 18636
rect 13236 18400 13321 18636
rect 13557 18400 13642 18636
rect 13878 18400 13963 18636
rect 14199 18400 14284 18636
rect 14520 18400 14605 18636
rect 14841 18400 15000 18636
rect 0 18300 15000 18400
rect 0 18064 143 18300
rect 379 18064 465 18300
rect 701 18064 787 18300
rect 1023 18064 1109 18300
rect 1345 18064 1431 18300
rect 1667 18064 1753 18300
rect 1989 18064 2075 18300
rect 2311 18064 2397 18300
rect 2633 18064 2719 18300
rect 2955 18064 3041 18300
rect 3277 18064 3363 18300
rect 3599 18064 3685 18300
rect 3921 18064 4007 18300
rect 4243 18064 4329 18300
rect 4565 18064 4651 18300
rect 4887 18064 4973 18300
rect 5209 18064 5295 18300
rect 5531 18064 9469 18300
rect 9705 18064 9790 18300
rect 10026 18064 10111 18300
rect 10347 18064 10432 18300
rect 10668 18064 10753 18300
rect 10989 18064 11074 18300
rect 11310 18064 11395 18300
rect 11631 18064 11716 18300
rect 11952 18064 12037 18300
rect 12273 18064 12358 18300
rect 12594 18064 12679 18300
rect 12915 18064 13000 18300
rect 13236 18064 13321 18300
rect 13557 18064 13642 18300
rect 13878 18064 13963 18300
rect 14199 18064 14284 18300
rect 14520 18064 14605 18300
rect 14841 18064 15000 18300
rect 0 17964 15000 18064
rect 0 17728 143 17964
rect 379 17728 465 17964
rect 701 17728 787 17964
rect 1023 17728 1109 17964
rect 1345 17728 1431 17964
rect 1667 17728 1753 17964
rect 1989 17728 2075 17964
rect 2311 17728 2397 17964
rect 2633 17728 2719 17964
rect 2955 17728 3041 17964
rect 3277 17728 3363 17964
rect 3599 17728 3685 17964
rect 3921 17728 4007 17964
rect 4243 17728 4329 17964
rect 4565 17728 4651 17964
rect 4887 17728 4973 17964
rect 5209 17728 5295 17964
rect 5531 17728 9469 17964
rect 9705 17728 9790 17964
rect 10026 17728 10111 17964
rect 10347 17728 10432 17964
rect 10668 17728 10753 17964
rect 10989 17728 11074 17964
rect 11310 17728 11395 17964
rect 11631 17728 11716 17964
rect 11952 17728 12037 17964
rect 12273 17728 12358 17964
rect 12594 17728 12679 17964
rect 12915 17728 13000 17964
rect 13236 17728 13321 17964
rect 13557 17728 13642 17964
rect 13878 17728 13963 17964
rect 14199 17728 14284 17964
rect 14520 17728 14605 17964
rect 14841 17728 15000 17964
rect 0 17628 15000 17728
rect 0 17392 143 17628
rect 379 17392 465 17628
rect 701 17392 787 17628
rect 1023 17392 1109 17628
rect 1345 17392 1431 17628
rect 1667 17392 1753 17628
rect 1989 17392 2075 17628
rect 2311 17392 2397 17628
rect 2633 17392 2719 17628
rect 2955 17392 3041 17628
rect 3277 17392 3363 17628
rect 3599 17392 3685 17628
rect 3921 17392 4007 17628
rect 4243 17392 4329 17628
rect 4565 17392 4651 17628
rect 4887 17392 4973 17628
rect 5209 17392 5295 17628
rect 5531 17392 9469 17628
rect 9705 17392 9790 17628
rect 10026 17392 10111 17628
rect 10347 17392 10432 17628
rect 10668 17392 10753 17628
rect 10989 17392 11074 17628
rect 11310 17392 11395 17628
rect 11631 17392 11716 17628
rect 11952 17392 12037 17628
rect 12273 17392 12358 17628
rect 12594 17392 12679 17628
rect 12915 17392 13000 17628
rect 13236 17392 13321 17628
rect 13557 17392 13642 17628
rect 13878 17392 13963 17628
rect 14199 17392 14284 17628
rect 14520 17392 14605 17628
rect 14841 17392 15000 17628
rect 0 17292 15000 17392
rect 0 17056 143 17292
rect 379 17056 465 17292
rect 701 17056 787 17292
rect 1023 17056 1109 17292
rect 1345 17056 1431 17292
rect 1667 17056 1753 17292
rect 1989 17056 2075 17292
rect 2311 17056 2397 17292
rect 2633 17056 2719 17292
rect 2955 17056 3041 17292
rect 3277 17056 3363 17292
rect 3599 17056 3685 17292
rect 3921 17056 4007 17292
rect 4243 17056 4329 17292
rect 4565 17056 4651 17292
rect 4887 17056 4973 17292
rect 5209 17056 5295 17292
rect 5531 17056 9469 17292
rect 9705 17056 9790 17292
rect 10026 17056 10111 17292
rect 10347 17056 10432 17292
rect 10668 17056 10753 17292
rect 10989 17056 11074 17292
rect 11310 17056 11395 17292
rect 11631 17056 11716 17292
rect 11952 17056 12037 17292
rect 12273 17056 12358 17292
rect 12594 17056 12679 17292
rect 12915 17056 13000 17292
rect 13236 17056 13321 17292
rect 13557 17056 13642 17292
rect 13878 17056 13963 17292
rect 14199 17056 14284 17292
rect 14520 17056 14605 17292
rect 14841 17056 15000 17292
rect 0 16956 15000 17056
rect 0 16720 143 16956
rect 379 16720 465 16956
rect 701 16720 787 16956
rect 1023 16720 1109 16956
rect 1345 16720 1431 16956
rect 1667 16720 1753 16956
rect 1989 16720 2075 16956
rect 2311 16720 2397 16956
rect 2633 16720 2719 16956
rect 2955 16720 3041 16956
rect 3277 16720 3363 16956
rect 3599 16720 3685 16956
rect 3921 16720 4007 16956
rect 4243 16720 4329 16956
rect 4565 16720 4651 16956
rect 4887 16720 4973 16956
rect 5209 16720 5295 16956
rect 5531 16720 9469 16956
rect 9705 16720 9790 16956
rect 10026 16720 10111 16956
rect 10347 16720 10432 16956
rect 10668 16720 10753 16956
rect 10989 16720 11074 16956
rect 11310 16720 11395 16956
rect 11631 16720 11716 16956
rect 11952 16720 12037 16956
rect 12273 16720 12358 16956
rect 12594 16720 12679 16956
rect 12915 16720 13000 16956
rect 13236 16720 13321 16956
rect 13557 16720 13642 16956
rect 13878 16720 13963 16956
rect 14199 16720 14284 16956
rect 14520 16720 14605 16956
rect 14841 16720 15000 16956
rect 0 16620 15000 16720
rect 0 16384 143 16620
rect 379 16384 465 16620
rect 701 16384 787 16620
rect 1023 16384 1109 16620
rect 1345 16384 1431 16620
rect 1667 16384 1753 16620
rect 1989 16384 2075 16620
rect 2311 16384 2397 16620
rect 2633 16384 2719 16620
rect 2955 16384 3041 16620
rect 3277 16384 3363 16620
rect 3599 16384 3685 16620
rect 3921 16384 4007 16620
rect 4243 16384 4329 16620
rect 4565 16384 4651 16620
rect 4887 16384 4973 16620
rect 5209 16384 5295 16620
rect 5531 16384 9469 16620
rect 9705 16384 9790 16620
rect 10026 16384 10111 16620
rect 10347 16384 10432 16620
rect 10668 16384 10753 16620
rect 10989 16384 11074 16620
rect 11310 16384 11395 16620
rect 11631 16384 11716 16620
rect 11952 16384 12037 16620
rect 12273 16384 12358 16620
rect 12594 16384 12679 16620
rect 12915 16384 13000 16620
rect 13236 16384 13321 16620
rect 13557 16384 13642 16620
rect 13878 16384 13963 16620
rect 14199 16384 14284 16620
rect 14520 16384 14605 16620
rect 14841 16384 15000 16620
rect 0 16284 15000 16384
rect 0 16048 143 16284
rect 379 16048 465 16284
rect 701 16048 787 16284
rect 1023 16048 1109 16284
rect 1345 16048 1431 16284
rect 1667 16048 1753 16284
rect 1989 16048 2075 16284
rect 2311 16048 2397 16284
rect 2633 16048 2719 16284
rect 2955 16048 3041 16284
rect 3277 16048 3363 16284
rect 3599 16048 3685 16284
rect 3921 16048 4007 16284
rect 4243 16048 4329 16284
rect 4565 16048 4651 16284
rect 4887 16048 4973 16284
rect 5209 16048 5295 16284
rect 5531 16048 9469 16284
rect 9705 16048 9790 16284
rect 10026 16048 10111 16284
rect 10347 16048 10432 16284
rect 10668 16048 10753 16284
rect 10989 16048 11074 16284
rect 11310 16048 11395 16284
rect 11631 16048 11716 16284
rect 11952 16048 12037 16284
rect 12273 16048 12358 16284
rect 12594 16048 12679 16284
rect 12915 16048 13000 16284
rect 13236 16048 13321 16284
rect 13557 16048 13642 16284
rect 13878 16048 13963 16284
rect 14199 16048 14284 16284
rect 14520 16048 14605 16284
rect 14841 16048 15000 16284
rect 0 15948 15000 16048
rect 0 15712 143 15948
rect 379 15712 465 15948
rect 701 15712 787 15948
rect 1023 15712 1109 15948
rect 1345 15712 1431 15948
rect 1667 15712 1753 15948
rect 1989 15712 2075 15948
rect 2311 15712 2397 15948
rect 2633 15712 2719 15948
rect 2955 15712 3041 15948
rect 3277 15712 3363 15948
rect 3599 15712 3685 15948
rect 3921 15712 4007 15948
rect 4243 15712 4329 15948
rect 4565 15712 4651 15948
rect 4887 15712 4973 15948
rect 5209 15712 5295 15948
rect 5531 15712 9469 15948
rect 9705 15712 9790 15948
rect 10026 15712 10111 15948
rect 10347 15712 10432 15948
rect 10668 15712 10753 15948
rect 10989 15712 11074 15948
rect 11310 15712 11395 15948
rect 11631 15712 11716 15948
rect 11952 15712 12037 15948
rect 12273 15712 12358 15948
rect 12594 15712 12679 15948
rect 12915 15712 13000 15948
rect 13236 15712 13321 15948
rect 13557 15712 13642 15948
rect 13878 15712 13963 15948
rect 14199 15712 14284 15948
rect 14520 15712 14605 15948
rect 14841 15712 15000 15948
rect 0 15612 15000 15712
rect 0 15376 143 15612
rect 379 15376 465 15612
rect 701 15376 787 15612
rect 1023 15376 1109 15612
rect 1345 15376 1431 15612
rect 1667 15376 1753 15612
rect 1989 15376 2075 15612
rect 2311 15376 2397 15612
rect 2633 15376 2719 15612
rect 2955 15376 3041 15612
rect 3277 15376 3363 15612
rect 3599 15376 3685 15612
rect 3921 15376 4007 15612
rect 4243 15376 4329 15612
rect 4565 15376 4651 15612
rect 4887 15376 4973 15612
rect 5209 15376 5295 15612
rect 5531 15376 9469 15612
rect 9705 15376 9790 15612
rect 10026 15376 10111 15612
rect 10347 15376 10432 15612
rect 10668 15376 10753 15612
rect 10989 15376 11074 15612
rect 11310 15376 11395 15612
rect 11631 15376 11716 15612
rect 11952 15376 12037 15612
rect 12273 15376 12358 15612
rect 12594 15376 12679 15612
rect 12915 15376 13000 15612
rect 13236 15376 13321 15612
rect 13557 15376 13642 15612
rect 13878 15376 13963 15612
rect 14199 15376 14284 15612
rect 14520 15376 14605 15612
rect 14841 15376 15000 15612
rect 0 15276 15000 15376
rect 0 15040 143 15276
rect 379 15040 465 15276
rect 701 15040 787 15276
rect 1023 15040 1109 15276
rect 1345 15040 1431 15276
rect 1667 15040 1753 15276
rect 1989 15040 2075 15276
rect 2311 15040 2397 15276
rect 2633 15040 2719 15276
rect 2955 15040 3041 15276
rect 3277 15040 3363 15276
rect 3599 15040 3685 15276
rect 3921 15040 4007 15276
rect 4243 15040 4329 15276
rect 4565 15040 4651 15276
rect 4887 15040 4973 15276
rect 5209 15040 5295 15276
rect 5531 15040 9469 15276
rect 9705 15040 9790 15276
rect 10026 15040 10111 15276
rect 10347 15040 10432 15276
rect 10668 15040 10753 15276
rect 10989 15040 11074 15276
rect 11310 15040 11395 15276
rect 11631 15040 11716 15276
rect 11952 15040 12037 15276
rect 12273 15040 12358 15276
rect 12594 15040 12679 15276
rect 12915 15040 13000 15276
rect 13236 15040 13321 15276
rect 13557 15040 13642 15276
rect 13878 15040 13963 15276
rect 14199 15040 14284 15276
rect 14520 15040 14605 15276
rect 14841 15040 15000 15276
rect 0 14940 15000 15040
rect 0 14704 143 14940
rect 379 14704 465 14940
rect 701 14704 787 14940
rect 1023 14704 1109 14940
rect 1345 14704 1431 14940
rect 1667 14704 1753 14940
rect 1989 14704 2075 14940
rect 2311 14704 2397 14940
rect 2633 14704 2719 14940
rect 2955 14704 3041 14940
rect 3277 14704 3363 14940
rect 3599 14704 3685 14940
rect 3921 14704 4007 14940
rect 4243 14704 4329 14940
rect 4565 14704 4651 14940
rect 4887 14704 4973 14940
rect 5209 14704 5295 14940
rect 5531 14704 9469 14940
rect 9705 14704 9790 14940
rect 10026 14704 10111 14940
rect 10347 14704 10432 14940
rect 10668 14704 10753 14940
rect 10989 14704 11074 14940
rect 11310 14704 11395 14940
rect 11631 14704 11716 14940
rect 11952 14704 12037 14940
rect 12273 14704 12358 14940
rect 12594 14704 12679 14940
rect 12915 14704 13000 14940
rect 13236 14704 13321 14940
rect 13557 14704 13642 14940
rect 13878 14704 13963 14940
rect 14199 14704 14284 14940
rect 14520 14704 14605 14940
rect 14841 14704 15000 14940
rect 0 14604 15000 14704
rect 0 14368 143 14604
rect 379 14368 465 14604
rect 701 14368 787 14604
rect 1023 14368 1109 14604
rect 1345 14368 1431 14604
rect 1667 14368 1753 14604
rect 1989 14368 2075 14604
rect 2311 14368 2397 14604
rect 2633 14368 2719 14604
rect 2955 14368 3041 14604
rect 3277 14368 3363 14604
rect 3599 14368 3685 14604
rect 3921 14368 4007 14604
rect 4243 14368 4329 14604
rect 4565 14368 4651 14604
rect 4887 14368 4973 14604
rect 5209 14368 5295 14604
rect 5531 14368 9469 14604
rect 9705 14368 9790 14604
rect 10026 14368 10111 14604
rect 10347 14368 10432 14604
rect 10668 14368 10753 14604
rect 10989 14368 11074 14604
rect 11310 14368 11395 14604
rect 11631 14368 11716 14604
rect 11952 14368 12037 14604
rect 12273 14368 12358 14604
rect 12594 14368 12679 14604
rect 12915 14368 13000 14604
rect 13236 14368 13321 14604
rect 13557 14368 13642 14604
rect 13878 14368 13963 14604
rect 14199 14368 14284 14604
rect 14520 14368 14605 14604
rect 14841 14368 15000 14604
rect 0 14268 15000 14368
rect 0 14032 143 14268
rect 379 14032 465 14268
rect 701 14032 787 14268
rect 1023 14032 1109 14268
rect 1345 14032 1431 14268
rect 1667 14032 1753 14268
rect 1989 14032 2075 14268
rect 2311 14032 2397 14268
rect 2633 14032 2719 14268
rect 2955 14032 3041 14268
rect 3277 14032 3363 14268
rect 3599 14032 3685 14268
rect 3921 14032 4007 14268
rect 4243 14032 4329 14268
rect 4565 14032 4651 14268
rect 4887 14032 4973 14268
rect 5209 14032 5295 14268
rect 5531 14032 9469 14268
rect 9705 14032 9790 14268
rect 10026 14032 10111 14268
rect 10347 14032 10432 14268
rect 10668 14032 10753 14268
rect 10989 14032 11074 14268
rect 11310 14032 11395 14268
rect 11631 14032 11716 14268
rect 11952 14032 12037 14268
rect 12273 14032 12358 14268
rect 12594 14032 12679 14268
rect 12915 14032 13000 14268
rect 13236 14032 13321 14268
rect 13557 14032 13642 14268
rect 13878 14032 13963 14268
rect 14199 14032 14284 14268
rect 14520 14032 14605 14268
rect 14841 14032 15000 14268
rect 0 14007 15000 14032
<< rm5 >>
tri 2404 34212 2424 34232 se
rect 2424 34212 12577 34232
tri 12577 34212 12597 34232 sw
tri 2389 34197 2404 34212 se
rect 2404 34197 2417 34212
tri 2417 34197 2432 34212 nw
tri 2361 34169 2389 34197 se
tri 2389 34169 2417 34197 nw
tri 12569 34184 12597 34212 ne
tri 12597 34184 12625 34212 sw
tri 2333 34141 2361 34169 se
tri 2361 34141 2389 34169 nw
tri 12597 34156 12625 34184 ne
tri 12625 34156 12653 34184 sw
tri 2305 34113 2333 34141 se
tri 2333 34113 2361 34141 nw
tri 12625 34128 12653 34156 ne
tri 12653 34128 12681 34156 sw
tri 2277 34085 2305 34113 se
tri 2305 34085 2333 34113 nw
tri 12653 34100 12681 34128 ne
tri 12681 34100 12709 34128 sw
tri 2249 34057 2277 34085 se
tri 2277 34057 2305 34085 nw
tri 12681 34072 12709 34100 ne
tri 12709 34072 12737 34100 sw
tri 2221 34029 2249 34057 se
tri 2249 34029 2277 34057 nw
tri 12709 34044 12737 34072 ne
tri 12737 34044 12765 34072 sw
tri 2193 34001 2221 34029 se
tri 2221 34001 2249 34029 nw
tri 12737 34016 12765 34044 ne
tri 12765 34016 12793 34044 sw
tri 2165 33973 2193 34001 se
tri 2193 33973 2221 34001 nw
tri 12765 33988 12793 34016 ne
tri 12793 33988 12821 34016 sw
tri 2137 33945 2165 33973 se
tri 2165 33945 2193 33973 nw
tri 12793 33960 12821 33988 ne
tri 12821 33960 12849 33988 sw
tri 2109 33917 2137 33945 se
tri 2137 33917 2165 33945 nw
tri 12821 33932 12849 33960 ne
tri 12849 33932 12877 33960 sw
tri 2081 33889 2109 33917 se
tri 2109 33889 2137 33917 nw
tri 12849 33904 12877 33932 ne
tri 12877 33904 12905 33932 sw
tri 2053 33861 2081 33889 se
tri 2081 33861 2109 33889 nw
tri 12877 33876 12905 33904 ne
tri 12905 33876 12933 33904 sw
tri 2025 33833 2053 33861 se
tri 2053 33833 2081 33861 nw
tri 12905 33848 12933 33876 ne
tri 12933 33848 12961 33876 sw
tri 1997 33805 2025 33833 se
tri 2025 33805 2053 33833 nw
tri 12933 33820 12961 33848 ne
tri 12961 33820 12989 33848 sw
tri 1969 33777 1997 33805 se
tri 1997 33777 2025 33805 nw
tri 12961 33792 12989 33820 ne
tri 12989 33792 13017 33820 sw
tri 1941 33749 1969 33777 se
tri 1969 33749 1997 33777 nw
tri 12989 33764 13017 33792 ne
tri 13017 33764 13045 33792 sw
tri 1913 33721 1941 33749 se
tri 1941 33721 1969 33749 nw
tri 13017 33736 13045 33764 ne
tri 13045 33736 13073 33764 sw
tri 1885 33693 1913 33721 se
tri 1913 33693 1941 33721 nw
tri 13045 33708 13073 33736 ne
tri 13073 33708 13101 33736 sw
tri 1857 33665 1885 33693 se
tri 1885 33665 1913 33693 nw
tri 13073 33680 13101 33708 ne
tri 13101 33680 13129 33708 sw
tri 1829 33637 1857 33665 se
tri 1857 33637 1885 33665 nw
tri 13101 33652 13129 33680 ne
tri 13129 33652 13157 33680 sw
tri 1801 33609 1829 33637 se
tri 1829 33609 1857 33637 nw
tri 13129 33624 13157 33652 ne
tri 13157 33624 13185 33652 sw
tri 1773 33581 1801 33609 se
tri 1801 33581 1829 33609 nw
tri 13157 33596 13185 33624 ne
tri 13185 33596 13213 33624 sw
tri 1745 33553 1773 33581 se
tri 1773 33553 1801 33581 nw
tri 13185 33568 13213 33596 ne
tri 13213 33568 13241 33596 sw
tri 1717 33525 1745 33553 se
tri 1745 33525 1773 33553 nw
tri 13213 33540 13241 33568 ne
tri 13241 33540 13269 33568 sw
tri 1689 33497 1717 33525 se
tri 1717 33497 1745 33525 nw
tri 13241 33512 13269 33540 ne
tri 13269 33512 13297 33540 sw
tri 1661 33469 1689 33497 se
tri 1689 33469 1717 33497 nw
tri 13269 33484 13297 33512 ne
tri 13297 33484 13325 33512 sw
tri 1633 33441 1661 33469 se
tri 1661 33441 1689 33469 nw
tri 13297 33456 13325 33484 ne
tri 13325 33456 13353 33484 sw
tri 1605 33413 1633 33441 se
tri 1633 33413 1661 33441 nw
tri 13325 33428 13353 33456 ne
tri 13353 33428 13381 33456 sw
tri 1577 33385 1605 33413 se
tri 1605 33385 1633 33413 nw
tri 13353 33400 13381 33428 ne
tri 13381 33400 13409 33428 sw
tri 1549 33357 1577 33385 se
tri 1577 33357 1605 33385 nw
tri 13381 33372 13409 33400 ne
tri 13409 33372 13437 33400 sw
tri 1521 33329 1549 33357 se
tri 1549 33329 1577 33357 nw
tri 13409 33344 13437 33372 ne
tri 13437 33344 13465 33372 sw
tri 1493 33301 1521 33329 se
tri 1521 33301 1549 33329 nw
tri 13437 33316 13465 33344 ne
tri 13465 33316 13493 33344 sw
tri 1465 33273 1493 33301 se
tri 1493 33273 1521 33301 nw
tri 13465 33288 13493 33316 ne
tri 13493 33288 13521 33316 sw
tri 1437 33245 1465 33273 se
tri 1465 33245 1493 33273 nw
tri 13493 33260 13521 33288 ne
tri 13521 33260 13549 33288 sw
tri 1409 33217 1437 33245 se
tri 1437 33217 1465 33245 nw
tri 13521 33232 13549 33260 ne
tri 13549 33232 13577 33260 sw
tri 1381 33189 1409 33217 se
tri 1409 33189 1437 33217 nw
tri 13549 33204 13577 33232 ne
tri 13577 33204 13605 33232 sw
tri 1353 33161 1381 33189 se
tri 1381 33161 1409 33189 nw
tri 13577 33178 13603 33204 ne
rect 13603 33186 13605 33204
tri 13605 33186 13623 33204 sw
tri 1333 33141 1353 33161 se
rect 1333 21069 1353 33141
tri 1353 33133 1381 33161 nw
tri 1333 21049 1353 21069 ne
tri 1353 21049 1381 21077 sw
tri 1353 21024 1378 21049 ne
rect 1378 21024 1381 21049
tri 1381 21024 1406 21049 sw
tri 1378 20996 1406 21024 ne
tri 1406 20996 1434 21024 sw
tri 1406 20968 1434 20996 ne
tri 1434 20968 1462 20996 sw
tri 13575 20994 13603 21022 se
rect 13603 21014 13623 33186
tri 13603 20994 13623 21014 nw
tri 1434 20940 1462 20968 ne
tri 1462 20940 1490 20968 sw
tri 13547 20966 13575 20994 se
tri 13575 20966 13603 20994 nw
tri 1462 20912 1490 20940 ne
tri 1490 20912 1518 20940 sw
tri 13519 20938 13547 20966 se
tri 13547 20938 13575 20966 nw
tri 1490 20884 1518 20912 ne
tri 1518 20884 1546 20912 sw
tri 13491 20910 13519 20938 se
tri 13519 20910 13547 20938 nw
tri 1518 20856 1546 20884 ne
tri 1546 20856 1574 20884 sw
tri 13463 20882 13491 20910 se
tri 13491 20882 13519 20910 nw
tri 1546 20828 1574 20856 ne
tri 1574 20828 1602 20856 sw
tri 13435 20854 13463 20882 se
tri 13463 20854 13491 20882 nw
tri 1574 20800 1602 20828 ne
tri 1602 20800 1630 20828 sw
tri 13407 20826 13435 20854 se
tri 13435 20826 13463 20854 nw
tri 1602 20772 1630 20800 ne
tri 1630 20772 1658 20800 sw
tri 13379 20798 13407 20826 se
tri 13407 20798 13435 20826 nw
tri 1630 20744 1658 20772 ne
tri 1658 20744 1686 20772 sw
tri 13351 20770 13379 20798 se
tri 13379 20770 13407 20798 nw
tri 1658 20716 1686 20744 ne
tri 1686 20716 1714 20744 sw
tri 13323 20742 13351 20770 se
tri 13351 20742 13379 20770 nw
tri 1686 20688 1714 20716 ne
tri 1714 20688 1742 20716 sw
tri 13295 20714 13323 20742 se
tri 13323 20714 13351 20742 nw
tri 1714 20660 1742 20688 ne
tri 1742 20660 1770 20688 sw
tri 13267 20686 13295 20714 se
tri 13295 20686 13323 20714 nw
tri 1742 20632 1770 20660 ne
tri 1770 20632 1798 20660 sw
tri 13239 20658 13267 20686 se
tri 13267 20658 13295 20686 nw
tri 1770 20604 1798 20632 ne
tri 1798 20604 1826 20632 sw
tri 13211 20630 13239 20658 se
tri 13239 20630 13267 20658 nw
tri 1798 20576 1826 20604 ne
tri 1826 20576 1854 20604 sw
tri 13183 20602 13211 20630 se
tri 13211 20602 13239 20630 nw
tri 1826 20548 1854 20576 ne
tri 1854 20548 1882 20576 sw
tri 13155 20574 13183 20602 se
tri 13183 20574 13211 20602 nw
tri 1854 20520 1882 20548 ne
tri 1882 20520 1910 20548 sw
tri 13127 20546 13155 20574 se
tri 13155 20546 13183 20574 nw
tri 1882 20492 1910 20520 ne
tri 1910 20492 1938 20520 sw
tri 13099 20518 13127 20546 se
tri 13127 20518 13155 20546 nw
tri 1910 20464 1938 20492 ne
tri 1938 20464 1966 20492 sw
tri 13071 20490 13099 20518 se
tri 13099 20490 13127 20518 nw
tri 1938 20436 1966 20464 ne
tri 1966 20436 1994 20464 sw
tri 13043 20462 13071 20490 se
tri 13071 20462 13099 20490 nw
tri 1966 20408 1994 20436 ne
tri 1994 20408 2022 20436 sw
tri 13015 20434 13043 20462 se
tri 13043 20434 13071 20462 nw
tri 1994 20380 2022 20408 ne
tri 2022 20380 2050 20408 sw
tri 12987 20406 13015 20434 se
tri 13015 20406 13043 20434 nw
tri 2022 20352 2050 20380 ne
tri 2050 20352 2078 20380 sw
tri 12959 20378 12987 20406 se
tri 12987 20378 13015 20406 nw
tri 2050 20324 2078 20352 ne
tri 2078 20324 2106 20352 sw
tri 12931 20350 12959 20378 se
tri 12959 20350 12987 20378 nw
tri 2078 20296 2106 20324 ne
tri 2106 20296 2134 20324 sw
tri 12903 20322 12931 20350 se
tri 12931 20322 12959 20350 nw
tri 2106 20268 2134 20296 ne
tri 2134 20268 2162 20296 sw
tri 12875 20294 12903 20322 se
tri 12903 20294 12931 20322 nw
tri 2134 20240 2162 20268 ne
tri 2162 20240 2190 20268 sw
tri 12847 20266 12875 20294 se
tri 12875 20266 12903 20294 nw
tri 2162 20212 2190 20240 ne
tri 2190 20212 2218 20240 sw
tri 12819 20238 12847 20266 se
tri 12847 20238 12875 20266 nw
tri 2190 20184 2218 20212 ne
tri 2218 20184 2246 20212 sw
tri 12791 20210 12819 20238 se
tri 12819 20210 12847 20238 nw
tri 2218 20156 2246 20184 ne
tri 2246 20156 2274 20184 sw
tri 12763 20182 12791 20210 se
tri 12791 20182 12819 20210 nw
tri 2246 20128 2274 20156 ne
tri 2274 20128 2302 20156 sw
tri 12735 20154 12763 20182 se
tri 12763 20154 12791 20182 nw
tri 2274 20100 2302 20128 ne
tri 2302 20100 2330 20128 sw
tri 12707 20126 12735 20154 se
tri 12735 20126 12763 20154 nw
tri 2302 20072 2330 20100 ne
tri 2330 20072 2358 20100 sw
tri 12679 20098 12707 20126 se
tri 12707 20098 12735 20126 nw
tri 2330 20044 2358 20072 ne
tri 2358 20044 2386 20072 sw
tri 12651 20070 12679 20098 se
tri 12679 20070 12707 20098 nw
tri 2358 20016 2386 20044 ne
tri 2386 20016 2414 20044 sw
tri 12623 20042 12651 20070 se
tri 12651 20042 12679 20070 nw
tri 2386 19988 2414 20016 ne
tri 2414 19988 2442 20016 sw
tri 12595 20014 12623 20042 se
tri 12623 20014 12651 20042 nw
tri 2414 19960 2442 19988 ne
tri 2442 19960 2470 19988 sw
tri 12567 19986 12595 20014 se
tri 12595 19986 12623 20014 nw
tri 2442 19932 2470 19960 ne
tri 2470 19932 2498 19960 sw
tri 12539 19958 12567 19986 se
tri 12567 19958 12595 19986 nw
tri 2470 19904 2498 19932 ne
tri 2498 19904 2526 19932 sw
tri 12511 19930 12539 19958 se
tri 12539 19930 12567 19958 nw
tri 12485 19904 12511 19930 se
rect 12511 19904 12513 19930
tri 12513 19904 12539 19930 nw
tri 2498 19884 2518 19904 ne
rect 2518 19884 12493 19904
tri 12493 19884 12513 19904 nw
<< glass >>
tri 1499 33090 2489 34080 se
rect 2489 33090 12509 34080
tri 12509 33090 13499 34080 sw
rect 1499 21070 13499 33090
tri 1499 20080 2489 21070 ne
rect 2489 20080 12509 21070
tri 12509 20080 13499 21070 nw
<< labels >>
flabel metal4 s 0 35157 254 40000 3 FreeSans 1015 0 0 0 VSSIO
port 4 nsew
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 1015 180 0 0 VSSIO
port 4 nsew
flabel metal4 s 6904 14009 8104 14209 0 FreeSans 1400 0 0 0 P_CORE
port 1 nsew
flabel metal5 s 2000 20574 12990 33596 0 FreeSans 3906 0 0 0 P_PAD
port 2 nsew
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 1015 180 0 0 VDDIO
port 3 nsew
flabel metal5 s 0 14007 254 18997 3 FreeSans 1015 0 0 0 VDDIO
port 3 nsew
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 1015 180 0 0 VDDIO
port 3 nsew
flabel metal4 s 0 14007 254 19000 3 FreeSans 1015 0 0 0 VDDIO
port 3 nsew
flabel metal5 s 0 35157 254 40000 3 FreeSans 1015 0 0 0 VSSIO
port 4 nsew
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 1015 180 0 0 VSSIO
port 4 nsew
flabel metal4 s 14873 37578 14873 37578 3 FreeSans 1015 180 0 0 VSSIO
flabel metal4 s 127 37578 127 37578 3 FreeSans 1015 0 0 0 VSSIO
flabel metal4 14746 35157 15000 40000 3 FreeSans 650 180 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_fd_io__com_bus_hookup_0.VSSIO
flabel metal4 14746 14007 15000 19000 3 FreeSans 650 180 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_fd_io__com_bus_hookup_0.VDDIO
flabel metal4 0 35157 254 40000 3 FreeSans 650 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_fd_io__com_bus_hookup_0.VSSIO
flabel metal4 0 14007 254 19000 3 FreeSans 650 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_fd_io__com_bus_hookup_0.VDDIO
flabel metal4 6904 14009 8104 14209 0 FreeSans 1400 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.P_CORE
flabel metal4 0 35157 254 40000 3 FreeSans 650 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VSSIO
flabel metal4 14746 35157 15000 40000 3 FreeSans 650 180 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VSSIO
flabel metal5 0 14007 254 18997 3 FreeSans 650 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VDDIO
flabel metal4 0 14007 254 19000 3 FreeSans 650 0 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VDDIO
flabel metal5 14746 14007 15000 18997 3 FreeSans 650 180 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VDDIO
flabel metal4 14746 14007 15000 19000 3 FreeSans 650 180 0 0 sky130_ef_io__minesd_pad_and_pg_0.sky130_ef_io__com_pg_esd_0.VDDIO
<< end >>
