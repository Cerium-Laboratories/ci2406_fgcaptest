magic
tech sky130A
magscale 1 2
timestamp 1717562480
<< xpolycontact >>
rect -35 19984 35 20416
rect -35 -20416 35 -19984
<< xpolyres >>
rect -35 -19984 35 19984
<< viali >>
rect -19 20001 19 20398
rect -19 -20398 19 -20001
<< metal1 >>
rect -25 20398 25 20410
rect -25 20001 -19 20398
rect 19 20001 25 20398
rect -25 19989 25 20001
rect -25 -20001 25 -19989
rect -25 -20398 -19 -20001
rect 19 -20398 25 -20001
rect -25 -20410 25 -20398
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 200 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 1.143meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
