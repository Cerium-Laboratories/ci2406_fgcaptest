magic
tech sky130A
timestamp 1717473404
<< nwell >>
rect -42 133 230 293
rect 357 133 1301 293
<< pwell >>
rect -14 -60 1273 55
<< mvnmos >>
rect 20 0 70 50
rect 99 0 149 50
rect 419 0 469 50
rect 498 0 548 50
rect 636 0 686 50
rect 715 0 765 50
rect 794 0 844 50
rect 873 0 923 50
rect 952 0 1002 50
rect 1031 0 1081 50
rect 1110 0 1160 50
rect 1189 0 1239 50
<< mvpmos >>
rect 20 166 70 216
rect 99 166 149 216
rect 419 166 469 216
rect 498 166 548 216
rect 636 166 686 216
rect 715 166 765 216
rect 794 166 844 216
rect 873 166 923 216
rect 952 166 1002 216
rect 1031 166 1081 216
rect 1110 166 1160 216
rect 1189 166 1239 216
<< mvndiff >>
rect -9 46 20 50
rect -9 4 -3 46
rect 14 4 20 46
rect -9 0 20 4
rect 70 46 99 50
rect 70 4 76 46
rect 93 4 99 46
rect 70 0 99 4
rect 149 46 178 50
rect 149 4 155 46
rect 172 4 178 46
rect 149 0 178 4
rect 390 46 419 50
rect 390 4 396 46
rect 413 4 419 46
rect 390 0 419 4
rect 469 46 498 50
rect 469 4 475 46
rect 492 4 498 46
rect 469 0 498 4
rect 548 46 577 50
rect 548 4 554 46
rect 571 4 577 46
rect 548 0 577 4
rect 607 46 636 50
rect 607 4 613 46
rect 630 4 636 46
rect 607 0 636 4
rect 686 46 715 50
rect 686 4 692 46
rect 709 4 715 46
rect 686 0 715 4
rect 765 46 794 50
rect 765 4 771 46
rect 788 4 794 46
rect 765 0 794 4
rect 844 46 873 50
rect 844 4 850 46
rect 867 4 873 46
rect 844 0 873 4
rect 923 46 952 50
rect 923 4 929 46
rect 946 4 952 46
rect 923 0 952 4
rect 1002 46 1031 50
rect 1002 4 1008 46
rect 1025 4 1031 46
rect 1002 0 1031 4
rect 1081 46 1110 50
rect 1081 4 1087 46
rect 1104 4 1110 46
rect 1081 0 1110 4
rect 1160 46 1189 50
rect 1160 4 1166 46
rect 1183 4 1189 46
rect 1160 0 1189 4
rect 1239 46 1268 50
rect 1239 4 1245 46
rect 1262 4 1268 46
rect 1239 0 1268 4
<< mvpdiff >>
rect -9 212 20 216
rect -9 170 -3 212
rect 14 170 20 212
rect -9 166 20 170
rect 70 212 99 216
rect 70 170 76 212
rect 93 170 99 212
rect 70 166 99 170
rect 149 212 178 216
rect 149 170 155 212
rect 172 170 178 212
rect 149 166 178 170
rect 390 212 419 216
rect 390 170 396 212
rect 413 170 419 212
rect 390 166 419 170
rect 469 212 498 216
rect 469 170 475 212
rect 492 170 498 212
rect 469 166 498 170
rect 548 212 577 216
rect 548 170 554 212
rect 571 170 577 212
rect 548 166 577 170
rect 607 212 636 216
rect 607 170 613 212
rect 630 170 636 212
rect 607 166 636 170
rect 686 212 715 216
rect 686 170 692 212
rect 709 170 715 212
rect 686 166 715 170
rect 765 212 794 216
rect 765 170 771 212
rect 788 170 794 212
rect 765 166 794 170
rect 844 212 873 216
rect 844 170 850 212
rect 867 170 873 212
rect 844 166 873 170
rect 923 212 952 216
rect 923 170 929 212
rect 946 170 952 212
rect 923 166 952 170
rect 1002 212 1031 216
rect 1002 170 1008 212
rect 1025 170 1031 212
rect 1002 166 1031 170
rect 1081 212 1110 216
rect 1081 170 1087 212
rect 1104 170 1110 212
rect 1081 166 1110 170
rect 1160 212 1189 216
rect 1160 170 1166 212
rect 1183 170 1189 212
rect 1160 166 1189 170
rect 1239 212 1268 216
rect 1239 170 1245 212
rect 1262 170 1268 212
rect 1239 166 1268 170
<< mvndiffc >>
rect -3 4 14 46
rect 76 4 93 46
rect 155 4 172 46
rect 396 4 413 46
rect 475 4 492 46
rect 554 4 571 46
rect 613 4 630 46
rect 692 4 709 46
rect 771 4 788 46
rect 850 4 867 46
rect 929 4 946 46
rect 1008 4 1025 46
rect 1087 4 1104 46
rect 1166 4 1183 46
rect 1245 4 1262 46
<< mvpdiffc >>
rect -3 170 14 212
rect 76 170 93 212
rect 155 170 172 212
rect 396 170 413 212
rect 475 170 492 212
rect 554 170 571 212
rect 613 170 630 212
rect 692 170 709 212
rect 771 170 788 212
rect 850 170 867 212
rect 929 170 946 212
rect 1008 170 1025 212
rect 1087 170 1104 212
rect 1166 170 1183 212
rect 1245 170 1262 212
<< mvpsubdiff >>
rect -3 -60 9 -43
rect 1250 -60 1262 -43
<< mvnsubdiff >>
rect -3 243 9 260
rect 185 243 197 260
rect 390 243 402 260
rect 1250 243 1262 260
<< mvpsubdiffcont >>
rect 9 -60 1250 -43
<< mvnsubdiffcont >>
rect 9 243 185 260
rect 402 243 1250 260
<< poly >>
rect 20 216 70 229
rect 99 216 149 229
rect 419 216 469 229
rect 498 216 548 229
rect 636 216 686 229
rect 715 216 765 229
rect 794 216 844 229
rect 873 216 923 229
rect 952 216 1002 229
rect 1031 216 1081 229
rect 1110 216 1160 229
rect 1189 216 1239 229
rect 20 140 70 166
rect 20 123 31 140
rect 59 123 70 140
rect 20 50 70 123
rect 99 97 149 166
rect 419 142 469 166
rect 419 125 430 142
rect 458 125 469 142
rect 419 120 469 125
rect 498 142 548 166
rect 498 125 509 142
rect 537 125 548 142
rect 498 120 548 125
rect 636 158 686 166
rect 715 158 765 166
rect 794 158 844 166
rect 873 158 923 166
rect 636 131 923 158
rect 99 80 110 97
rect 138 80 149 97
rect 636 114 647 131
rect 675 114 923 131
rect 636 112 923 114
rect 952 158 1002 166
rect 1031 158 1081 166
rect 1110 158 1160 166
rect 1189 158 1239 166
rect 952 141 1239 158
rect 99 50 149 80
rect 419 91 469 96
rect 419 74 430 91
rect 458 74 469 91
rect 419 50 469 74
rect 498 91 548 96
rect 498 74 509 91
rect 537 74 548 91
rect 498 50 548 74
rect 636 58 765 112
rect 636 50 686 58
rect 715 50 765 58
rect 794 86 923 91
rect 794 69 810 86
rect 827 69 923 86
rect 794 58 923 69
rect 794 50 844 58
rect 873 50 923 58
rect 952 75 957 141
rect 991 112 1239 141
rect 991 75 1081 112
rect 952 58 1081 75
rect 952 50 1002 58
rect 1031 50 1081 58
rect 1110 86 1239 91
rect 1110 69 1126 86
rect 1143 69 1239 86
rect 1110 58 1239 69
rect 1110 50 1160 58
rect 1189 50 1239 58
rect 20 -13 70 0
rect 99 -13 149 0
rect 419 -13 469 0
rect 498 -13 548 0
rect 636 -13 686 0
rect 715 -13 765 0
rect 794 -13 844 0
rect 873 -13 923 0
rect 952 -13 1002 0
rect 1031 -13 1081 0
rect 1110 -13 1160 0
rect 1189 -13 1239 0
<< polycont >>
rect 31 123 59 140
rect 430 125 458 142
rect 509 125 537 142
rect 110 80 138 97
rect 647 114 675 131
rect 430 74 458 91
rect 509 74 537 91
rect 810 69 827 86
rect 957 75 991 141
rect 1126 69 1143 86
<< locali >>
rect -3 254 9 260
rect 185 254 197 260
rect -3 243 3 254
rect 191 243 197 254
rect 390 254 402 260
rect 1250 254 1262 260
rect 390 243 396 254
rect -3 212 14 220
rect -3 97 14 170
rect 76 212 93 220
rect 76 162 93 170
rect 155 212 172 220
rect 31 140 59 148
rect 31 115 59 123
rect -3 46 14 80
rect 110 97 138 105
rect 110 72 138 80
rect 155 57 172 170
rect -3 -4 14 4
rect 76 46 93 54
rect 76 -21 93 4
rect 155 -4 172 4
rect 396 212 413 220
rect 475 212 492 237
rect 475 162 492 170
rect 554 212 571 220
rect 396 46 413 159
rect 430 142 458 150
rect 430 117 458 125
rect 509 148 514 165
rect 532 148 537 165
rect 509 142 537 148
rect 509 117 537 125
rect 554 139 571 170
rect 613 212 630 237
rect 613 162 630 170
rect 692 212 709 220
rect 692 162 709 170
rect 771 212 788 237
rect 771 162 788 170
rect 850 212 867 220
rect 850 162 867 170
rect 929 212 946 237
rect 929 162 946 170
rect 1008 212 1025 220
rect 957 141 991 149
rect 554 131 675 139
rect 571 114 647 131
rect 554 106 675 114
rect 430 91 458 99
rect 430 66 458 74
rect 509 91 537 99
rect 509 66 537 74
rect 396 -4 413 4
rect 475 46 492 54
rect 475 -21 492 4
rect 554 46 571 106
rect 771 69 810 86
rect 827 69 867 86
rect 771 54 867 69
rect 957 67 991 75
rect 1087 212 1104 237
rect 1087 162 1104 170
rect 1166 212 1183 220
rect 1166 162 1183 170
rect 1245 212 1262 237
rect 1245 162 1262 170
rect 554 -4 571 4
rect 613 46 630 54
rect 613 -21 630 4
rect 692 46 709 54
rect 692 -4 709 4
rect 771 46 788 54
rect 771 -4 788 4
rect 850 46 867 54
rect 850 -4 867 4
rect 929 46 946 54
rect 929 -4 946 4
rect 1008 46 1025 132
rect 1008 -4 1025 4
rect 1087 69 1126 86
rect 1143 69 1183 86
rect 1087 54 1183 69
rect 1087 46 1104 54
rect 1087 -4 1104 4
rect 1166 46 1183 54
rect 1166 -4 1183 4
rect 1245 46 1262 54
rect 1245 -4 1262 4
rect 771 -21 946 -4
rect 1087 -21 1262 -4
rect -3 -43 1262 -38
rect -3 -60 9 -43
rect 1250 -60 1262 -43
<< viali >>
rect 3 243 9 254
rect 9 243 185 254
rect 185 243 191 254
rect 396 243 402 254
rect 402 243 1250 254
rect 1250 243 1262 254
rect 3 237 191 243
rect 396 237 1262 243
rect 76 170 93 212
rect 36 123 54 140
rect -3 80 14 97
rect 115 80 133 97
rect 155 46 172 57
rect 155 40 172 46
rect 396 170 413 176
rect 396 159 413 170
rect 435 125 453 142
rect 514 148 532 165
rect 692 170 709 212
rect 850 170 867 212
rect 1008 170 1025 212
rect 554 114 571 131
rect 652 114 670 131
rect 435 74 453 91
rect 514 74 532 91
rect 954 75 957 109
rect 957 75 988 109
rect 1008 132 1025 170
rect 1166 170 1183 212
rect 692 4 709 46
rect -3 -38 1262 -21
<< metal1 >>
rect -3 254 197 257
rect -3 237 3 254
rect 191 237 197 254
rect -3 234 197 237
rect 390 254 1268 257
rect 390 237 396 254
rect 1262 237 1268 254
rect 390 234 1268 237
rect 73 212 96 234
rect 692 215 709 218
rect 850 215 867 218
rect 73 170 76 212
rect 93 170 96 212
rect 689 212 712 215
rect 73 164 96 170
rect 393 176 538 182
rect 393 159 396 176
rect 413 165 538 176
rect 689 170 692 212
rect 709 170 712 212
rect 689 167 712 170
rect 847 212 870 215
rect 847 170 850 212
rect 867 170 870 212
rect 847 167 870 170
rect 1005 212 1028 218
rect 1166 215 1183 218
rect 413 159 514 165
rect 393 153 416 159
rect 508 148 514 159
rect 532 148 538 165
rect 30 140 60 148
rect 508 145 538 148
rect 30 123 36 140
rect 54 123 60 140
rect 30 115 60 123
rect 429 142 494 145
rect 429 125 435 142
rect 453 131 494 142
rect 551 134 574 137
rect 551 131 676 134
rect 453 125 554 131
rect 429 122 554 125
rect 473 114 554 122
rect 571 114 652 131
rect 670 114 676 131
rect 551 111 676 114
rect 692 112 709 167
rect 850 112 867 167
rect 1005 132 1008 212
rect 1025 166 1028 212
rect 1163 212 1186 215
rect 1163 170 1166 212
rect 1183 170 1186 212
rect 1163 166 1186 170
rect 1025 132 1301 166
rect 1005 129 1301 132
rect 1008 126 1301 129
rect 551 108 574 111
rect 692 109 1301 112
rect -6 100 17 103
rect -6 97 459 100
rect -6 80 -3 97
rect 14 80 115 97
rect 133 91 459 97
rect 133 80 435 91
rect -6 77 435 80
rect -6 74 17 77
rect 429 74 435 77
rect 453 74 459 91
rect 429 71 459 74
rect 508 91 538 94
rect 508 74 514 91
rect 532 74 538 91
rect 152 57 175 63
rect 508 57 538 74
rect 152 40 155 57
rect 172 40 538 57
rect 692 78 954 109
rect 692 72 810 78
rect 827 75 954 78
rect 988 75 1301 109
rect 827 72 1301 75
rect 692 49 709 72
rect 152 34 538 40
rect 689 46 712 49
rect 689 4 692 46
rect 709 4 712 46
rect 689 1 712 4
rect 692 -2 709 1
rect -9 -21 1268 -18
rect -9 -38 -3 -21
rect 1262 -38 1268 -21
rect -9 -41 1268 -38
<< labels >>
flabel metal1 30 115 60 148 0 FreeSans 160 0 0 0 in
port 1 nsew
flabel locali -3 122 14 139 0 FreeSans 80 90 0 0 in_b
flabel locali 155 116 172 143 0 FreeSans 80 90 0 0 in_bb
flabel metal1 73 234 96 257 0 FreeSans 160 0 0 0 vdd_l
port 4 nsew
flabel metal1 -9 -41 14 -18 0 FreeSans 160 0 0 0 vss
port 6 nsew
flabel metal1 1261 72 1301 112 0 FreeSans 160 0 0 0 out
port 3 nsew
flabel metal1 1261 126 1301 166 0 FreeSans 160 0 0 0 out_b
port 2 nsew
flabel locali 554 80 571 97 0 FreeSans 80 0 0 0 t1
flabel locali 396 116 413 133 0 FreeSans 80 0 0 0 t2
flabel metal1 1245 234 1268 257 0 FreeSans 160 0 0 0 vdd_h
port 5 nsew
<< end >>
