magic
tech sky130A
magscale 1 2
timestamp 1717155884
<< error_s >>
rect 838 -1496 1300 -1336
rect 838 -2662 1300 -2502
<< nwell >>
rect 2410 -2164 3204 -1834
rect 6436 -2010 7910 -1988
<< mvnsubdiff >>
rect 6436 -2010 7910 -1988
<< polycont >>
rect 1138 -1449 1202 -1387
rect 1138 -2612 1204 -2550
<< locali >>
rect 1122 -1378 1218 -1371
rect 1122 -1456 1132 -1378
rect 1210 -1456 1218 -1378
rect 1122 -1465 1218 -1456
rect 1122 -2543 1220 -2534
rect 1122 -2621 1132 -2543
rect 1210 -2621 1220 -2543
rect 1122 -2628 1220 -2621
<< viali >>
rect 1132 -1387 1210 -1378
rect 1132 -1449 1138 -1387
rect 1138 -1449 1202 -1387
rect 1202 -1449 1210 -1387
rect 1132 -1456 1210 -1449
rect 1132 -2550 1210 -2543
rect 1132 -2612 1138 -2550
rect 1138 -2612 1204 -2550
rect 1204 -2612 1210 -2550
rect 1132 -2621 1210 -2612
<< metal1 >>
rect 1126 -1372 1216 -1366
rect 1120 -1462 1126 -1372
rect 1216 -1462 1222 -1372
rect 1126 -1468 1216 -1462
rect 6328 -2016 7872 -1982
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via1 >>
rect 1126 -1378 1216 -1372
rect 1126 -1456 1132 -1378
rect 1132 -1456 1210 -1378
rect 1210 -1456 1216 -1378
rect 1126 -1462 1216 -1456
rect 1126 -2543 1216 -2537
rect 1126 -2621 1132 -2543
rect 1132 -2621 1210 -2543
rect 1210 -2621 1216 -2543
rect 1126 -2627 1216 -2621
<< metal2 >>
rect 1126 -1372 1216 -1366
rect 1122 -1457 1126 -1377
rect 1216 -1457 1220 -1377
rect 1126 -1468 1216 -1462
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via2 >>
rect 1131 -1457 1211 -1377
rect 1131 -2622 1211 -2542
<< metal3 >>
rect 1126 -1377 1216 -1366
rect 1126 -1457 1131 -1377
rect 1211 -1457 1216 -1377
rect 1126 -1870 1216 -1457
rect 152 -2128 2208 -1870
rect 1126 -2538 1216 -2532
rect 1121 -2542 1221 -2538
rect 1121 -2622 1131 -2542
rect 1211 -2622 1221 -2542
rect 1121 -2626 1221 -2622
rect 1126 -2632 1216 -2626
<< mimcap >>
rect 180 -2008 2180 -1898
rect 180 -2078 1136 -2008
rect 1206 -2078 2180 -2008
rect 180 -2100 2180 -2078
<< mimcapcontact >>
rect 1136 -2078 1206 -2008
<< metal4 >>
rect 1126 -2008 1216 -1998
rect 1126 -2078 1136 -2008
rect 1206 -2078 1216 -2008
rect 1126 -2632 1216 -2078
use fgcell_amp  fgcell_amp_0
timestamp 1717155884
transform 1 0 0 0 -1 -6798
box 140 -5818 7976 -4698
use fgcell_amp  fgcell_amp_1
timestamp 1717155884
transform 1 0 0 0 1 2800
box 140 -5818 7976 -4698
<< end >>
