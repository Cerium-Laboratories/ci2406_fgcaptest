** sch_path: /Users/dalejulson/Desktop/OpenCircuitDesign/ci2406_fgcaptest/xschem/fgcell_MiM_cap_1_1.sch
**.subckt fgcell_MiM_cap_1_1 vinj vinj_en_b vtun vctrl vsrc
*.ipin vinj
*.ipin vinj_en_b
*.ipin vtun
*.ipin vctrl
*.ipin vsrc
x1 vinj vinj_en_b net1 vtun vctrl vsrc GND fgcell
XC1 net1 GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**** begin user architecture code
.lib /Users/dalejulson/Desktop/OpenCircuitDesign/open_pdks/sky130//sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  fgcell.sym # of pins=7
** sym_path: /Users/dalejulson/Desktop/OpenCircuitDesign/ci2406_fgcaptest/xschem/fgcell.sym
** sch_path: /Users/dalejulson/Desktop/OpenCircuitDesign/ci2406_fgcaptest/xschem/fgcell.sch
.subckt fgcell vinj vinj_en_b vfg vtun vctrl vsrc VGND
*.ipin vctrl
*.ipin vtun
*.ipin vinj
*.ipin vinj_en_b
*.ipin vsrc
*.opin vfg
*.ipin VGND
XC1 vfg vtun vtun sky130_fd_pr__cap_var_hvt W=0.5 L=0.5 VM=1 m=1
XM1 vsrc vfg net1 vinj sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 vinj_en_b vinj vinj sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vctrl vfg vctrl vctrl sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
