magic
tech sky130A
timestamp 1717160680
<< error_p >>
rect 349 14374 580 14454
rect 2349 14374 2580 14454
rect 4349 14374 4580 14454
rect 6349 14374 6580 14454
rect 8349 14374 8580 14454
rect 10349 14374 10580 14454
rect 12349 14374 12580 14454
rect 14349 14374 14580 14454
rect 16349 14374 16580 14454
rect 18349 14374 18580 14454
rect 349 12874 580 12954
rect 2349 12874 2580 12954
rect 4349 12874 4580 12954
rect 6349 12874 6580 12954
rect 8349 12874 8580 12954
rect 10349 12874 10580 12954
rect 12349 12874 12580 12954
rect 14349 12874 14580 12954
rect 16349 12874 16580 12954
rect 18349 12874 18580 12954
rect 349 11374 580 11454
rect 2349 11374 2580 11454
rect 4349 11374 4580 11454
rect 6349 11374 6580 11454
rect 8349 11374 8580 11454
rect 10349 11374 10580 11454
rect 12349 11374 12580 11454
rect 14349 11374 14580 11454
rect 16349 11374 16580 11454
rect 18349 11374 18580 11454
rect 349 9874 580 9954
rect 2349 9874 2580 9954
rect 4349 9874 4580 9954
rect 6349 9874 6580 9954
rect 8349 9874 8580 9954
rect 10349 9874 10580 9954
rect 12349 9874 12580 9954
rect 14349 9874 14580 9954
rect 16349 9874 16580 9954
rect 18349 9874 18580 9954
rect 349 8374 580 8454
rect 2349 8374 2580 8454
rect 4349 8374 4580 8454
rect 6349 8374 6580 8454
rect 8349 8374 8580 8454
rect 10349 8374 10580 8454
rect 12349 8374 12580 8454
rect 14349 8374 14580 8454
rect 16349 8374 16580 8454
rect 18349 8374 18580 8454
rect 349 6874 580 6954
rect 2349 6874 2580 6954
rect 4349 6874 4580 6954
rect 6349 6874 6580 6954
rect 8349 6874 8580 6954
rect 10349 6874 10580 6954
rect 12349 6874 12580 6954
rect 14349 6874 14580 6954
rect 16349 6874 16580 6954
rect 18349 6874 18580 6954
rect 349 5374 580 5454
rect 2349 5374 2580 5454
rect 4349 5374 4580 5454
rect 6349 5374 6580 5454
rect 8349 5374 8580 5454
rect 10349 5374 10580 5454
rect 12349 5374 12580 5454
rect 14349 5374 14580 5454
rect 16349 5374 16580 5454
rect 18349 5374 18580 5454
rect 349 3874 580 3954
rect 2349 3874 2580 3954
rect 4349 3874 4580 3954
rect 6349 3874 6580 3954
rect 8349 3874 8580 3954
rect 10349 3874 10580 3954
rect 12349 3874 12580 3954
rect 14349 3874 14580 3954
rect 16349 3874 16580 3954
rect 18349 3874 18580 3954
rect 349 2374 580 2454
rect 2349 2374 2580 2454
rect 4349 2374 4580 2454
rect 6349 2374 6580 2454
rect 8349 2374 8580 2454
rect 10349 2374 10580 2454
rect 12349 2374 12580 2454
rect 14349 2374 14580 2454
rect 16349 2374 16580 2454
rect 18349 2374 18580 2454
rect 349 874 580 954
rect 2349 874 2580 954
rect 4349 874 4580 954
rect 6349 874 6580 954
rect 8349 874 8580 954
rect 10349 874 10580 954
rect 12349 874 12580 954
rect 14349 874 14580 954
rect 16349 874 16580 954
rect 18349 874 18580 954
use fgcell_amp  fgcell_amp_0
array 0 9 2000 0 9 1500
timestamp 1717158785
transform 1 0 -70 0 1 3605
box 70 -3605 2053 -2482
<< end >>
