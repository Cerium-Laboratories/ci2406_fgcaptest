magic
tech sky130A
magscale 1 2
timestamp 1717349067
<< nwell >>
rect 3204 -1834 3668 -1804
rect 2410 -2164 3668 -1834
rect 3204 -2194 3668 -2164
<< polycont >>
rect 1142 -1445 1200 -1387
rect 1140 -2612 1202 -2548
<< locali >>
rect 1126 -1378 1216 -1371
rect 1126 -1456 1132 -1378
rect 1210 -1456 1216 -1378
rect 1126 -1461 1216 -1456
rect 1124 -2543 1218 -2532
rect 1124 -2621 1132 -2543
rect 1210 -2621 1218 -2543
rect 1124 -2628 1218 -2621
<< viali >>
rect 1132 -1387 1210 -1378
rect 1132 -1445 1142 -1387
rect 1142 -1445 1200 -1387
rect 1200 -1445 1210 -1387
rect 1132 -1456 1210 -1445
rect 1132 -2548 1210 -2543
rect 1132 -2612 1140 -2548
rect 1140 -2612 1202 -2548
rect 1202 -2612 1210 -2548
rect 1132 -2621 1210 -2612
<< metal1 >>
rect 1126 -1372 1216 -1366
rect 1120 -1462 1126 -1372
rect 1216 -1462 1222 -1372
rect 1126 -1468 1216 -1462
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via1 >>
rect 1126 -1378 1216 -1372
rect 1126 -1456 1132 -1378
rect 1132 -1456 1210 -1378
rect 1210 -1456 1216 -1378
rect 1126 -1462 1216 -1456
rect 1126 -2543 1216 -2537
rect 1126 -2621 1132 -2543
rect 1132 -2621 1210 -2543
rect 1210 -2621 1216 -2543
rect 1126 -2627 1216 -2621
<< metal2 >>
rect 1126 -1372 1216 -1366
rect 1122 -1457 1126 -1377
rect 1216 -1457 1220 -1377
rect 1126 -1468 1216 -1462
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via2 >>
rect 1131 -1457 1211 -1377
rect 1131 -2622 1211 -2542
<< metal3 >>
rect 1126 -1377 1216 -1366
rect 1126 -1457 1131 -1377
rect 1211 -1457 1216 -1377
rect 1126 -1874 1216 -1457
rect 1086 -2134 1356 -1874
rect 1126 -2538 1216 -2532
rect 1121 -2626 1127 -2538
rect 1215 -2626 1221 -2538
rect 1126 -2632 1216 -2626
<< via3 >>
rect 1127 -2542 1215 -2538
rect 1127 -2622 1131 -2542
rect 1131 -2622 1211 -2542
rect 1211 -2622 1215 -2542
rect 1127 -2626 1215 -2622
<< mimcap >>
rect 1116 -2014 1316 -1904
rect 1116 -2084 1136 -2014
rect 1206 -2084 1316 -2014
rect 1116 -2104 1316 -2084
<< mimcapcontact >>
rect 1136 -2084 1206 -2014
<< metal4 >>
rect 1126 -2014 1216 -2004
rect 1126 -2084 1136 -2014
rect 1206 -2084 1216 -2014
rect 1126 -2538 1216 -2084
rect 1126 -2626 1127 -2538
rect 1215 -2626 1216 -2538
rect 1126 -2632 1216 -2626
use fgcell_amp  fgcell_amp_0
timestamp 1717349067
transform 1 0 0 0 -1 -6798
box 140 -7210 4106 -4964
use fgcell_amp  fgcell_amp_1
timestamp 1717349067
transform 1 0 0 0 1 2800
box 140 -7210 4106 -4964
<< end >>
