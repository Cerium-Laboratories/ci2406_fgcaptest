magic
tech sky130A
timestamp 1717191602
<< nwell >>
rect 10 860 570 1450
<< pwell >>
rect 40 -10 540 760
<< mvnmos >>
rect 100 600 200 750
rect 250 600 350 750
rect 100 300 200 450
rect 250 300 350 450
rect 100 0 200 150
rect 250 0 350 150
<< mvpmos >>
rect 100 1200 200 1350
rect 250 1200 350 1350
rect 100 900 200 1050
rect 250 900 350 1050
<< mvndiff >>
rect 50 740 100 750
rect 50 610 60 740
rect 90 610 100 740
rect 50 600 100 610
rect 200 740 250 750
rect 200 610 210 740
rect 240 610 250 740
rect 200 600 250 610
rect 350 740 400 750
rect 350 610 360 740
rect 390 610 400 740
rect 350 600 400 610
rect 50 440 100 450
rect 50 310 60 440
rect 90 310 100 440
rect 50 300 100 310
rect 200 300 250 450
rect 350 440 400 450
rect 350 310 360 440
rect 390 310 400 440
rect 350 300 400 310
rect 50 140 100 150
rect 50 10 60 140
rect 90 10 100 140
rect 50 0 100 10
rect 200 140 250 150
rect 200 10 210 140
rect 240 10 250 140
rect 200 0 250 10
rect 350 140 400 150
rect 350 10 360 140
rect 390 10 400 140
rect 350 0 400 10
<< mvpdiff >>
rect 50 1340 100 1350
rect 50 1210 60 1340
rect 90 1210 100 1340
rect 50 1200 100 1210
rect 200 1340 250 1350
rect 200 1210 210 1340
rect 240 1210 250 1340
rect 200 1200 250 1210
rect 350 1340 400 1350
rect 350 1210 360 1340
rect 390 1210 400 1340
rect 350 1200 400 1210
rect 50 1040 100 1050
rect 50 910 60 1040
rect 90 910 100 1040
rect 50 900 100 910
rect 200 1040 250 1050
rect 200 910 210 1040
rect 240 910 250 1040
rect 200 900 250 910
rect 350 1040 400 1050
rect 350 910 360 1040
rect 390 910 400 1040
rect 350 900 400 910
<< mvndiffc >>
rect 60 610 90 740
rect 210 610 240 740
rect 360 610 390 740
rect 60 310 90 440
rect 360 310 390 440
rect 60 10 90 140
rect 210 10 240 140
rect 360 10 390 140
<< mvpdiffc >>
rect 60 1210 90 1340
rect 210 1210 240 1340
rect 360 1210 390 1340
rect 60 910 90 1040
rect 210 910 240 1040
rect 360 910 390 1040
<< mvpsubdiff >>
rect 470 480 530 500
rect 470 120 490 480
rect 510 120 530 480
rect 470 110 530 120
<< mvnsubdiff >>
rect 470 1340 530 1350
rect 470 1100 490 1340
rect 510 1100 530 1340
rect 470 1090 530 1100
<< mvpsubdiffcont >>
rect 490 120 510 480
<< mvnsubdiffcont >>
rect 490 1100 510 1340
<< poly >>
rect 100 1350 200 1370
rect 250 1350 350 1370
rect 100 1180 200 1200
rect 250 1180 350 1200
rect 100 1170 350 1180
rect 100 1150 260 1170
rect 340 1150 350 1170
rect 100 1140 350 1150
rect 100 1050 200 1070
rect 250 1050 350 1070
rect 100 880 200 900
rect 250 880 350 900
rect 100 870 350 880
rect 100 850 110 870
rect 190 850 350 870
rect 100 840 350 850
rect 100 750 200 770
rect 250 750 350 770
rect 100 590 200 600
rect 250 590 350 600
rect 100 580 350 590
rect 100 540 110 580
rect 190 540 350 580
rect 100 530 350 540
rect 100 450 200 470
rect 250 450 350 470
rect 100 290 200 300
rect 250 290 350 300
rect 100 280 350 290
rect 100 260 260 280
rect 340 260 350 280
rect 100 250 350 260
rect 100 150 200 170
rect 250 150 350 170
rect 100 -70 200 0
rect 250 -30 350 0
rect 250 -50 260 -30
rect 340 -50 350 -30
rect 250 -70 350 -50
<< polycont >>
rect 260 1150 340 1170
rect 110 850 190 870
rect 110 540 190 580
rect 260 260 340 280
rect 260 -50 340 -30
<< locali >>
rect 60 1340 90 1350
rect 60 1200 90 1210
rect 210 1340 240 1350
rect 10 1040 90 1050
rect 10 910 13 1040
rect 37 910 60 1040
rect 10 900 90 910
rect 210 1040 240 1210
rect 360 1340 400 1350
rect 390 1210 400 1340
rect 360 1180 400 1210
rect 260 1170 400 1180
rect 340 1150 400 1170
rect 260 1130 400 1150
rect 490 1340 510 1350
rect 490 1090 510 1100
rect 210 900 240 910
rect 360 1040 390 1050
rect 360 900 390 910
rect 60 880 90 900
rect 60 870 200 880
rect 60 850 110 870
rect 190 850 200 870
rect 60 840 200 850
rect 60 740 90 750
rect 60 580 90 610
rect 210 740 240 750
rect 210 600 240 610
rect 360 740 390 750
rect 360 600 390 610
rect 60 540 110 580
rect 190 540 200 580
rect 360 517 530 520
rect 360 473 366 517
rect 407 480 530 517
rect 407 473 490 480
rect 50 440 100 450
rect 50 310 60 440
rect 90 310 100 440
rect 50 220 100 310
rect 360 440 490 473
rect 390 310 490 440
rect 360 300 490 310
rect 260 280 340 290
rect 260 250 340 260
rect 50 170 250 220
rect 10 140 90 150
rect 10 10 60 140
rect 10 0 90 10
rect 200 140 250 170
rect 200 10 210 140
rect 240 10 250 140
rect 200 0 250 10
rect 360 140 390 150
rect 470 120 490 300
rect 510 120 530 480
rect 470 110 530 120
rect 360 0 390 10
rect 260 -30 340 -20
rect 260 -60 340 -50
<< viali >>
rect 63 1210 87 1340
rect 13 910 37 1040
rect 363 1210 387 1340
rect 490 1100 510 1340
rect 210 910 240 1040
rect 363 910 387 1040
rect 63 610 87 740
rect 210 610 240 740
rect 363 610 387 740
rect 366 473 407 517
rect 260 260 340 280
rect 63 10 87 140
rect 363 10 387 140
rect 490 120 510 480
rect 260 -50 340 -30
<< metal1 >>
rect 200 1380 520 1430
rect 60 1340 90 1350
rect 60 1210 63 1340
rect 87 1210 90 1340
rect 10 1040 40 1050
rect 10 910 13 1040
rect 37 910 40 1040
rect 10 150 40 910
rect 60 740 90 1210
rect 200 1040 250 1380
rect 360 1340 460 1350
rect 360 1210 363 1340
rect 387 1210 460 1340
rect 360 1200 460 1210
rect 200 910 210 1040
rect 240 910 250 1040
rect 200 900 250 910
rect 360 1040 390 1050
rect 360 910 363 1040
rect 387 910 390 1040
rect 360 900 390 910
rect 360 750 361 900
rect 387 750 390 900
rect 60 610 63 740
rect 87 610 90 740
rect 60 600 90 610
rect 200 740 250 750
rect 200 610 210 740
rect 240 610 250 740
rect 200 520 250 610
rect 360 740 390 750
rect 360 610 363 740
rect 387 610 390 740
rect 360 600 390 610
rect 200 517 413 520
rect 200 480 366 517
rect 360 473 366 480
rect 407 473 413 517
rect 360 470 413 473
rect 250 290 350 300
rect 250 260 260 290
rect 340 260 350 290
rect 250 250 350 260
rect 430 150 460 1200
rect 480 1340 520 1380
rect 480 1100 490 1340
rect 510 1100 520 1340
rect 480 1090 520 1100
rect 10 140 90 150
rect 10 10 63 140
rect 87 10 90 140
rect 10 0 90 10
rect 360 140 460 150
rect 360 10 363 140
rect 387 10 460 140
rect 480 480 530 490
rect 480 120 490 480
rect 510 120 530 480
rect 480 100 530 120
rect 360 0 460 10
rect 250 -30 350 -20
rect 250 -60 260 -30
rect 340 -60 350 -30
rect 250 -70 350 -60
<< via1 >>
rect 361 750 387 900
rect 260 280 340 290
rect 260 260 340 280
rect 260 -50 340 -30
rect 260 -60 340 -50
<< metal2 >>
rect 358 900 390 903
rect 358 750 361 900
rect 387 750 390 900
rect 358 747 390 750
rect 250 290 350 300
rect 250 260 260 290
rect 340 260 350 290
rect 250 250 350 260
rect 250 -30 350 -20
rect 250 -60 260 -30
rect 340 -60 350 -30
rect 250 -70 350 -60
<< labels >>
flabel metal1 480 100 530 150 0 FreeSans 80 0 0 0 VSS
port 3 nsew ground default
flabel metal1 200 1380 250 1430 0 FreeSans 80 0 0 0 VDD
port 4 nsew
flabel poly 100 -70 200 -20 0 FreeSans 80 0 0 0 v1
port 1 nsew analog input
flabel metal2 250 -70 350 -20 0 FreeSans 80 0 0 0 v2
port 2 nsew analog input
flabel metal1 60 1090 90 1120 0 FreeSans 160 0 0 0 int2
flabel metal1 10 780 40 810 0 FreeSans 160 0 0 0 int4
flabel mvndiff 200 300 250 450 0 FreeSans 160 0 0 0 int5
flabel metal2 358 747 390 903 0 FreeSans 160 0 0 0 vout
port 6 nsew
flabel pwell 470 510 520 560 0 FreeSans 160 0 0 0 VSS
flabel metal2 250 250 350 300 0 FreeSans 80 0 0 0 vb
port 5 nsew analog input
flabel metal1 430 1090 460 1120 0 FreeSans 160 0 0 0 int3
flabel locali 50 170 100 220 0 FreeSans 160 0 0 0 int1
<< end >>
