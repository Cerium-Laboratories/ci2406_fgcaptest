* NGSPICE file created from top_fgcaptest.ext - technology: sky130A

.subckt pad_minesd_short P_PAD P_CORE VDDIO VSSIO
R0 P_CORE P_PAD sky130_fd_pr__res_generic_m5 w=252.96 l=0.1
X0 P_CORE VDDIO sky130_fd_pr__diode_pd2nw_11v0 perim=1.02e+08 area=5e+13
X1 VSSIO P_CORE sky130_fd_pr__diode_pw2nd_11v0 perim=1.02e+08 area=5e+13
**devattr s=7137360,22068 d=7137360,22068
.ends

.subckt vtun_pad pad sky130_ef_io__bare_pad_0/VSUBS sky130_ef_io__bare_pad_0/PAD GND
X0 sky130_ef_io__bare_pad_0/PAD GND sky130_ef_io__bare_pad_0/VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=728.88
X1 a_5600_9600# sky130_ef_io__bare_pad_0/PAD sky130_fd_pr__res_generic_po w=7 l=24
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt array_column_decode a[3] a[2] a[1] a[0] w[15] w[14] w[13] w[12] w[11] w[10]
+ w[9] w[7] w[6] w[5] w[4] w[3] w[2] w[1] w[0] w[8] VGND VPWR
Xx3 a[2] VGND VGND VPWR VPWR x3/Y sky130_fd_sc_hd__inv_1
Xx2 a[3] VGND VGND VPWR VPWR x2/Y sky130_fd_sc_hd__inv_1
Xx4 a[1] VGND VGND VPWR VPWR x6/B sky130_fd_sc_hd__inv_1
Xx5 a[0] VGND VGND VPWR VPWR x8/A sky130_fd_sc_hd__inv_1
Xx6 x8/A x6/B VGND VGND VPWR VPWR x6/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand2_2_0 a[0] x6/B VGND VGND VPWR VPWR sky130_fd_sc_hd__nand2_2_0/Y
+ sky130_fd_sc_hd__nand2_2
Xx8 x8/A a[1] VGND VGND VPWR VPWR x8/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_1[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xx9 a[0] a[1] VGND VGND VPWR VPWR x9/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xx10 x3/Y x2/Y VGND VGND VPWR VPWR x10/Y sky130_fd_sc_hd__nand2_2
Xx11 a[2] x2/Y VGND VGND VPWR VPWR x11/Y sky130_fd_sc_hd__nand2_2
Xx12 x3/Y a[3] VGND VGND VPWR VPWR x12/Y sky130_fd_sc_hd__nand2_2
Xx13 a[2] a[3] VGND VGND VPWR VPWR x13/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nor3_1_0[0] x8/Y x13/Y VGND VGND VGND VPWR VPWR w[14] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[1] x6/Y x13/Y VGND VGND VGND VPWR VPWR w[12] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[2] x8/Y x12/Y VGND VGND VGND VPWR VPWR w[10] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[3] x6/Y x12/Y VGND VGND VGND VPWR VPWR w[8] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[4] x8/Y x11/Y VGND VGND VGND VPWR VPWR w[6] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[5] x6/Y x11/Y VGND VGND VGND VPWR VPWR w[4] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[6] x8/Y x10/Y VGND VGND VGND VPWR VPWR w[2] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[7] x6/Y x10/Y VGND VGND VGND VPWR VPWR w[0] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[0] x9/Y x13/Y VGND VGND VGND VPWR VPWR w[15] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[1] sky130_fd_sc_hd__nand2_2_0/Y x13/Y VGND VGND VGND VPWR
+ VPWR w[13] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[2] x9/Y x12/Y VGND VGND VGND VPWR VPWR w[11] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[3] sky130_fd_sc_hd__nand2_2_0/Y x12/Y VGND VGND VGND VPWR
+ VPWR w[9] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[4] x9/Y x11/Y VGND VGND VGND VPWR VPWR w[7] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[5] sky130_fd_sc_hd__nand2_2_0/Y x11/Y VGND VGND VGND VPWR
+ VPWR w[5] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[6] x9/Y x10/Y VGND VGND VGND VPWR VPWR w[3] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[7] sky130_fd_sc_hd__nand2_2_0/Y x10/Y VGND VGND VGND VPWR
+ VPWR w[1] sky130_fd_sc_hd__nor3_1
.ends

.subckt fgcell vinj vinj_en_b vtun vctrl vsrc VGND vfg
X0 a_697_110# vfg vsrc vinj sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 vfg vtun VGND sky130_fd_pr__cap_var w=1 l=0.5
X2 vinj vinj_en_b a_697_110# vinj sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X3 vctrl vfg vctrl vctrl sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.58 ps=5.16 w=1 l=0.5
.ends

.subckt diffamp_nmos v1 v2 VSS VDD vb vout
X0 int3 int3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X1 int1 v1 int4 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X2 int5 vb int1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X3 VSS int2 int2 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X4 VSS vb int5 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X5 VDD int4 int4 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X6 vout int2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X7 VDD int3 int2 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.375 pd=2 as=0.75 ps=4 w=1.5 l=1
X8 int3 v2 int1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
X9 vout int4 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=4 as=0.375 ps=2 w=1.5 l=1
.ends

.subckt tg5v0 vin vout en en_b vdd vss
X0 vout en vin vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 vout en vin vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 vin en vout vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X3 vin en vout vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X4 vout en vin vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X5 vout en_b vin vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X6 vout en_b vin vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X7 vin en vout vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X8 vin en vout vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X9 vin en_b vout vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X10 vin en_b vout vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X11 vout en vin vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X12 vout en_b vin vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X13 vin en_b vout vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X14 vin en_b vout vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X15 vout en_b vin vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt fgcell_amp_MOS_cap_thin_poly tg5v0_0/vout vdd vtun x1/vctrl row_en vsrc row_en_b
+ VGND x2/vb x1/vinj
Xx1 x1/vinj row_en_b vtun x1/vctrl vsrc VGND x2/v1 fgcell
Xx2 x2/v1 x2/v2 VGND vdd x2/vb x2/v2 diffamp_nmos
Xtg5v0_0 x2/v2 tg5v0_0/vout row_en row_en_b x1/vinj VGND tg5v0
X0 a_1282_n6014# x2/v1 a_1282_n6014# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=4.275 pd=34.58 as=4.275 ps=34.58 w=8.01 l=0.5
.ends

.subckt fgcell_amp_MOS_cap_thick_poly vout vdd row_en_b x1/vtun VSRC x1/vctrl row_en
+ VGND x2/vb vinj
Xx1 vinj row_en_b x1/vtun x1/vctrl VSRC VGND x2/v1 fgcell
Xx2 x2/v1 x2/v2 VGND vdd x2/vb x2/v2 diffamp_nmos
Xtg5v0_0 x2/v2 vout row_en row_en_b vinj VGND tg5v0
.ends

.subckt array_core_block5 fgcell_amp_MOS_cap_thick_poly_0[3|6]/vout fgcell_amp_MOS_cap_thin_poly_0[0|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|5]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/VSRC fgcell_amp_MOS_cap_thin_poly_0[0|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|5]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|6]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[1|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[2|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[4|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[3|1]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/row_en fgcell_amp_MOS_cap_thin_poly_0[3|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|3]/vsrc fgcell_amp_MOS_cap_thick_poly_0[2|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/vdd fgcell_amp_MOS_cap_thick_poly_0[2|3]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/vsrc fgcell_amp_MOS_cap_thick_poly_0[1|6]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/vinj fgcell_amp_MOS_cap_thin_poly_0[1|7]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/vout fgcell_amp_MOS_cap_thick_poly_0[0|7]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[4|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|2]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|9]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/vout fgcell_amp_MOS_cap_thick_poly_0[2|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|7]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/vdd fgcell_amp_MOS_cap_thick_poly_0[4|8]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[0|2]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|1]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[4|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[3|8]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|3]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[4|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/row_en fgcell_amp_MOS_cap_thick_poly_0[3|9]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[1|8]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[4|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|9]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[0|1]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/vsrc fgcell_amp_MOS_cap_thick_poly_0[3|6]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|5]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/vout fgcell_amp_MOS_cap_thin_poly_0[0|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|7]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|3]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|0]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/vtun fgcell_amp_MOS_cap_thin_poly_0[3|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/vsrc fgcell_amp_MOS_cap_thick_poly_0[4|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|6]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/vout fgcell_amp_MOS_cap_thin_poly_0[3|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/vtun fgcell_amp_MOS_cap_thin_poly_0[0|1]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/vinj fgcell_amp_MOS_cap_thin_poly_0[1|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/vout fgcell_amp_MOS_cap_thin_poly_0[3|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|6]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|8]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/vout fgcell_amp_MOS_cap_thin_poly_0[3|0]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[3|0]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[3|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/VSRC fgcell_amp_MOS_cap_thin_poly_0[0|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[3|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[4|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|5]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|7]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[0|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|4]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/vinj fgcell_amp_MOS_cap_thin_poly_0[4|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[2|8]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[3|4]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|8]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|3]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|6]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|5]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|8]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/vtun fgcell_amp_MOS_cap_thick_poly_0[2|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/vtun fgcell_amp_MOS_cap_thin_poly_0[3|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[4|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|6]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/vout fgcell_amp_MOS_cap_thin_poly_0[0|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[2|0]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[3|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/VSRC fgcell_amp_MOS_cap_thin_poly_0[3|3]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|8]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[0|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[0|2]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|6]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[2|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|8]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[4|2]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/VSRC fgcell_amp_MOS_cap_thin_poly_0[1|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/vtun fgcell_amp_MOS_cap_thick_poly_0[4|1]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|7]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[2|1]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|4]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[0|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/vout fgcell_amp_MOS_cap_thick_poly_0[1|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[4|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/vsrc fgcell_amp_MOS_cap_thick_poly_0[2|5]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/row_en fgcell_amp_MOS_cap_thin_poly_0[1|8]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/vout fgcell_amp_MOS_cap_thick_poly_0[1|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/vinj fgcell_amp_MOS_cap_thin_poly_0[3|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|6]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/vinj fgcell_amp_MOS_cap_thin_poly_0[2|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[2|3]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[2|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/vtun fgcell_amp_MOS_cap_thick_poly_0[2|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|0]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[4|3]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|9]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/vtun fgcell_amp_MOS_cap_thin_poly_0[2|2]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[3|8]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|6]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/vinj fgcell_amp_MOS_cap_thin_poly_0[1|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[3|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/VSRC fgcell_amp_MOS_cap_thin_poly_0[0|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/vinj fgcell_amp_MOS_cap_thick_poly_0[0|5]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[2|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|0]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/vout fgcell_amp_MOS_cap_thick_poly_0[1|1]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|2]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|4]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/vtun fgcell_amp_MOS_cap_thick_poly_0[3|3]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|2]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|7]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[0|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/vout fgcell_amp_MOS_cap_thin_poly_0[1|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|2]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/vinj fgcell_amp_MOS_cap_thin_poly_0[2|8]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/row_en fgcell_amp_MOS_cap_thick_poly_0[0|3]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/vtun fgcell_amp_MOS_cap_thin_poly_0[0|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|7]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|5]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[1|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/vtun fgcell_amp_MOS_cap_thick_poly_0[2|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[2|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/vsrc fgcell_amp_MOS_cap_thick_poly_0[0|6]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|8]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|9]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|9]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|4]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|0]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|0]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[3|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/vtun fgcell_amp_MOS_cap_thin_poly_0[3|5]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[2|3]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|0]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|0]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/vout fgcell_amp_MOS_cap_thin_poly_0[0|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[4|4]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|1]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/VSRC fgcell_amp_MOS_cap_thin_poly_0[1|1]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|0]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/VSRC fgcell_amp_MOS_cap_thin_poly_0[0|8]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/vout fgcell_amp_MOS_cap_thin_poly_0[3|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|6]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[2|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|6]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|1]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/vout fgcell_amp_MOS_cap_thick_poly_0[4|3]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|7]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[2|1]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/vtun fgcell_amp_MOS_cap_thick_poly_0[0|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[2|2]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[4|5]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/vout fgcell_amp_MOS_cap_thick_poly_0[3|2]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[0|0]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/vdd fgcell_amp_MOS_cap_thick_poly_0[2|2]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/vsrc fgcell_amp_MOS_cap_thick_poly_0[2|9]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[3|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|1]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[2|4]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/vtun fgcell_amp_MOS_cap_thin_poly_0[2|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[0|6]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|4]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/vinj fgcell_amp_MOS_cap_thick_poly_0[1|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/vsrc fgcell_amp_MOS_cap_thick_poly_0[0|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|8]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|4]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/vdd fgcell_amp_MOS_cap_thick_poly_0[4|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/vinj fgcell_amp_MOS_cap_thin_poly_0[4|7]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|3]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/vtun fgcell_amp_MOS_cap_thin_poly_0[2|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/vout fgcell_amp_MOS_cap_thick_poly_0[2|8]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/vtun fgcell_amp_MOS_cap_thick_poly_0[2|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[0|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[4|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|9]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|4]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|9]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|0]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[2|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|0]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[1|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|6]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|3]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[4|7]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/vout fgcell_amp_MOS_cap_thin_poly_0[2|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[0|4]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|1]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|2]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|8]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|4]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/vinj fgcell_amp_MOS_cap_thin_poly_0[0|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[0|2]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/vinj fgcell_amp_MOS_cap_thin_poly_0[3|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|1]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/vinj fgcell_amp_MOS_cap_thin_poly_0[1|0]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|9]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[3|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|4]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|9]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|8]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/vinj fgcell_amp_MOS_cap_thick_poly_0[4|8]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|9]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|8]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/vtun fgcell_amp_MOS_cap_thin_poly_0[4|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/vinj fgcell_amp_MOS_cap_thick_poly_0[0|9]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|9]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/vinj fgcell_amp_MOS_cap_thin_poly_0[3|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/vtun fgcell_amp_MOS_cap_thick_poly_0[0|0]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|8]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/VSRC fgcell_amp_MOS_cap_thin_poly_0[4|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/row_en fgcell_amp_MOS_cap_thick_poly_0[4|3]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/vtun fgcell_amp_MOS_cap_thin_poly_0[4|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|9]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|1]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|0]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[2|7]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/vout fgcell_amp_MOS_cap_thin_poly_0[0|9]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|8]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|7]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|1]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[3|9]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|5]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/row_en fgcell_amp_MOS_cap_thick_poly_0[4|7]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[2|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/VSRC fgcell_amp_MOS_cap_thin_poly_0[3|3]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|8]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|1]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[2|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[3|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|9]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[1|2]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[3|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|7]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/vsrc fgcell_amp_MOS_cap_thick_poly_0[0|5]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/vinj fgcell_amp_MOS_cap_thick_poly_0[0|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/VSRC fgcell_amp_MOS_cap_thin_poly_0[2|9]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|4]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|3]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|4]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/vsrc fgcell_amp_MOS_cap_thick_poly_0[0|6]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|8]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/vinj fgcell_amp_MOS_cap_thin_poly_0[2|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/vsrc fgcell_amp_MOS_cap_thick_poly_0[4|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/row_en fgcell_amp_MOS_cap_thick_poly_0[3|0]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/vinj fgcell_amp_MOS_cap_thick_poly_0[2|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|7]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|9]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/vtun fgcell_amp_MOS_cap_thick_poly_0[4|6]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|9]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[4|0]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[2|1]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/VSRC fgcell_amp_MOS_cap_thin_poly_0[3|8]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|2]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|1]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[2|2]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|2]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|4]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/vout fgcell_amp_MOS_cap_thick_poly_0[4|5]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[3|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[2|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[1|8]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[4|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|4]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[4|3]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/vdd fgcell_amp_MOS_cap_thick_poly_0[2|5]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[2|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[1|1]/VSRC
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/row_en fgcell_amp_MOS_cap_thick_poly_0[1|3]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/vdd fgcell_amp_MOS_cap_thick_poly_0[4|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[0|8]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[2|2]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/vout fgcell_amp_MOS_cap_thick_poly_0[0|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[4|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[3|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|5]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/row_en fgcell_amp_MOS_cap_thick_poly_0[4|6]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|0]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|9]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[2|4]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/vinj fgcell_amp_MOS_cap_thin_poly_0[0|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|6]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/x1/vctrl fgcell_amp_MOS_cap_thick_poly_0[0|8]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|3]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/vinj fgcell_amp_MOS_cap_thick_poly_0[3|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/vtun fgcell_amp_MOS_cap_thin_poly_0[1|3]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/vinj fgcell_amp_MOS_cap_thin_poly_0[4|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/vtun fgcell_amp_MOS_cap_thin_poly_0[4|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|5]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|1]/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/vinj fgcell_amp_MOS_cap_thick_poly_0[3|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|3]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/row_en fgcell_amp_MOS_cap_thin_poly_0[3|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|8]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/VSRC fgcell_amp_MOS_cap_thin_poly_0[0|9]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/vtun fgcell_amp_MOS_cap_thin_poly_0[2|0]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|9]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|8]/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/vtun fgcell_amp_MOS_cap_thick_poly_0[3|0]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|2]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/vinj fgcell_amp_MOS_cap_thin_poly_0[3|5]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[3|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[1|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|4]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/row_en fgcell_amp_MOS_cap_thick_poly_0[2|1]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|2]/x1/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[4|9]/vout
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/x2/vb fgcell_amp_MOS_cap_thick_poly_0[1|8]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[0|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/row_en fgcell_amp_MOS_cap_thin_poly_0[2|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[2|3]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/x1/vtun fgcell_amp_MOS_cap_thick_poly_0[2|8]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[3|7]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[1|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[0|5]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|9]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[0|2]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|5]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|2]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[4|9]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|7]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|7]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/vdd fgcell_amp_MOS_cap_thick_poly_0[3|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[4|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/vdd fgcell_amp_MOS_cap_thick_poly_0[0|4]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/vinj fgcell_amp_MOS_cap_thin_poly_0[3|6]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/x1/vinj fgcell_amp_MOS_cap_thin_poly_0[3|9]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/row_en fgcell_amp_MOS_cap_thin_poly_0[1|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/x1/vinj fgcell_amp_MOS_cap_thick_poly_0[0|4]/x1/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|8]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/x1/vtun fgcell_amp_MOS_cap_thin_poly_0[4|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|5]/vsrc
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/vinj fgcell_amp_MOS_cap_thick_poly_0[4|1]/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/vsrc fgcell_amp_MOS_cap_thick_poly_0[0|2]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/vtun fgcell_amp_MOS_cap_thin_poly_0[1|8]/row_en_b
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/vinj fgcell_amp_MOS_cap_thin_poly_0[0|3]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|7]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/tg5v0_0/vout fgcell_amp_MOS_cap_thin_poly_0[0|5]/vdd
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|3]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/vout fgcell_amp_MOS_cap_thin_poly_0[0|6]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/row_en fgcell_amp_MOS_cap_thin_poly_0[3|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/vsrc fgcell_amp_MOS_cap_thick_poly_0[2|3]/vinj
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/vdd fgcell_amp_MOS_cap_thick_poly_0[1|2]/row_en
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/vinj fgcell_amp_MOS_cap_thin_poly_0[0|7]/vsrc
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|3]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/row_en fgcell_amp_MOS_cap_thin_poly_0[0|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/row_en fgcell_amp_MOS_cap_thin_poly_0[4|4]/x2/vb
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/vtun fgcell_amp_MOS_cap_thick_poly_0[0|1]/vinj
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|9]/vtun fgcell_amp_MOS_cap_thick_poly_0[1|5]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/tg5v0_0/vout fgcell_amp_MOS_cap_thick_poly_0[4|5]/row_en_b
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/row_en fgcell_amp_MOS_cap_thick_poly_0[4|4]/VSRC
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/row_en_b fgcell_amp_MOS_cap_thin_poly_0[4|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/vsrc fgcell_amp_MOS_cap_thick_poly_0[1|3]/row_en
Xfgcell_amp_MOS_cap_thin_poly_0[0|0] fgcell_amp_MOS_cap_thin_poly_0[0|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|0]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|0] fgcell_amp_MOS_cap_thin_poly_0[1|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|0]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|0] fgcell_amp_MOS_cap_thin_poly_0[2|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|0]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|0] fgcell_amp_MOS_cap_thin_poly_0[3|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|0]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|0] fgcell_amp_MOS_cap_thin_poly_0[4|0]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|0]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|0]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|0]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|0]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|0]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|0]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|1] fgcell_amp_MOS_cap_thin_poly_0[0|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|1]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|1]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|1] fgcell_amp_MOS_cap_thin_poly_0[1|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|1]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|1]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|1] fgcell_amp_MOS_cap_thin_poly_0[2|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|1]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|1]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|1] fgcell_amp_MOS_cap_thin_poly_0[3|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|1]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|1]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|1] fgcell_amp_MOS_cap_thin_poly_0[4|1]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|1]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|1]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|1]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|1]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|1]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|1]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|2] fgcell_amp_MOS_cap_thin_poly_0[0|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|2]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|2]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|2] fgcell_amp_MOS_cap_thin_poly_0[1|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|2]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|2]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|2] fgcell_amp_MOS_cap_thin_poly_0[2|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|2]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|2]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|2] fgcell_amp_MOS_cap_thin_poly_0[3|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|2]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|2]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|2] fgcell_amp_MOS_cap_thin_poly_0[4|2]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|2]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|2]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|2]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|2]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|2]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|2]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|3] fgcell_amp_MOS_cap_thin_poly_0[0|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|3]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|3]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|3] fgcell_amp_MOS_cap_thin_poly_0[1|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|3]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|3]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|3] fgcell_amp_MOS_cap_thin_poly_0[2|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|3]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|3]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|3] fgcell_amp_MOS_cap_thin_poly_0[3|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|3]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|3]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|3] fgcell_amp_MOS_cap_thin_poly_0[4|3]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|3]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|3]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|3]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|3]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|3]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|3]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|4] fgcell_amp_MOS_cap_thin_poly_0[0|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|4]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|4]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|4] fgcell_amp_MOS_cap_thin_poly_0[1|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|4]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|4]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|4] fgcell_amp_MOS_cap_thin_poly_0[2|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|4]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|4]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|4] fgcell_amp_MOS_cap_thin_poly_0[3|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|4]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|4]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|4] fgcell_amp_MOS_cap_thin_poly_0[4|4]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|4]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|4]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|4]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|4]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|4]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|4]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|4]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|4]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|5] fgcell_amp_MOS_cap_thin_poly_0[0|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|5]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|5] fgcell_amp_MOS_cap_thin_poly_0[1|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|5]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|5] fgcell_amp_MOS_cap_thin_poly_0[2|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|5]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|5] fgcell_amp_MOS_cap_thin_poly_0[3|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|5]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|5] fgcell_amp_MOS_cap_thin_poly_0[4|5]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|5]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|5]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|5]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|5]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|5]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|5]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|6] fgcell_amp_MOS_cap_thin_poly_0[0|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|6]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|6]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|6] fgcell_amp_MOS_cap_thin_poly_0[1|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|6]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|6]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|6] fgcell_amp_MOS_cap_thin_poly_0[2|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|6]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|6]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|6] fgcell_amp_MOS_cap_thin_poly_0[3|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|6]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|6]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|6] fgcell_amp_MOS_cap_thin_poly_0[4|6]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|6]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|6]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|6]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|6]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|6]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|6]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|7] fgcell_amp_MOS_cap_thin_poly_0[0|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|7]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|7]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|7] fgcell_amp_MOS_cap_thin_poly_0[1|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|7]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|7]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|7] fgcell_amp_MOS_cap_thin_poly_0[2|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|7]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|7]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|7] fgcell_amp_MOS_cap_thin_poly_0[3|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|7]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|7]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|7] fgcell_amp_MOS_cap_thin_poly_0[4|7]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|7]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|7]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|7]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|7]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|7]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|7]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|7]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|7]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|8] fgcell_amp_MOS_cap_thin_poly_0[0|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|8]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|8]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|8] fgcell_amp_MOS_cap_thin_poly_0[1|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|8]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|8]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|8] fgcell_amp_MOS_cap_thin_poly_0[2|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|8]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|8]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|8] fgcell_amp_MOS_cap_thin_poly_0[3|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|8]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|8]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|8] fgcell_amp_MOS_cap_thin_poly_0[4|8]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|8]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|8]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|8]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|8]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|8]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|8]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[0|9] fgcell_amp_MOS_cap_thin_poly_0[0|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[0|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[0|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[0|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[0|9]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[0|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[0|9]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[1|9] fgcell_amp_MOS_cap_thin_poly_0[1|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[1|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[1|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[1|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[1|9]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[1|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[1|9]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[2|9] fgcell_amp_MOS_cap_thin_poly_0[2|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[2|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[2|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[2|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[2|9]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[2|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[2|9]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[3|9] fgcell_amp_MOS_cap_thin_poly_0[3|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[3|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[3|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[3|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[3|9]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[3|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[3|9]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thin_poly_0[4|9] fgcell_amp_MOS_cap_thin_poly_0[4|9]/tg5v0_0/vout
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/vdd fgcell_amp_MOS_cap_thin_poly_0[4|9]/vtun
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/x1/vctrl fgcell_amp_MOS_cap_thin_poly_0[4|9]/row_en
+ fgcell_amp_MOS_cap_thin_poly_0[4|9]/vsrc fgcell_amp_MOS_cap_thin_poly_0[4|9]/row_en_b
+ VSUBS fgcell_amp_MOS_cap_thin_poly_0[4|9]/x2/vb fgcell_amp_MOS_cap_thin_poly_0[4|9]/x1/vinj
+ fgcell_amp_MOS_cap_thin_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|0] fgcell_amp_MOS_cap_thick_poly_0[0|0]/vout fgcell_amp_MOS_cap_thick_poly_0[0|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|0]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|0] fgcell_amp_MOS_cap_thick_poly_0[1|0]/vout fgcell_amp_MOS_cap_thick_poly_0[1|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|0]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|0] fgcell_amp_MOS_cap_thick_poly_0[2|0]/vout fgcell_amp_MOS_cap_thick_poly_0[2|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|0]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|0] fgcell_amp_MOS_cap_thick_poly_0[3|0]/vout fgcell_amp_MOS_cap_thick_poly_0[3|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|0]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|0] fgcell_amp_MOS_cap_thick_poly_0[4|0]/vout fgcell_amp_MOS_cap_thick_poly_0[4|0]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|0]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|0]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|0]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|0]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|1] fgcell_amp_MOS_cap_thick_poly_0[0|1]/vout fgcell_amp_MOS_cap_thick_poly_0[0|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|1]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|1] fgcell_amp_MOS_cap_thick_poly_0[1|1]/vout fgcell_amp_MOS_cap_thick_poly_0[1|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|1]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|1] fgcell_amp_MOS_cap_thick_poly_0[2|1]/vout fgcell_amp_MOS_cap_thick_poly_0[2|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|1]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|1] fgcell_amp_MOS_cap_thick_poly_0[3|1]/vout fgcell_amp_MOS_cap_thick_poly_0[3|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|1]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|1] fgcell_amp_MOS_cap_thick_poly_0[4|1]/vout fgcell_amp_MOS_cap_thick_poly_0[4|1]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|1]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|1]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|1]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|1]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|2] fgcell_amp_MOS_cap_thick_poly_0[0|2]/vout fgcell_amp_MOS_cap_thick_poly_0[0|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|2]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|2] fgcell_amp_MOS_cap_thick_poly_0[1|2]/vout fgcell_amp_MOS_cap_thick_poly_0[1|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|2]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|2] fgcell_amp_MOS_cap_thick_poly_0[2|2]/vout fgcell_amp_MOS_cap_thick_poly_0[2|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|2]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|2] fgcell_amp_MOS_cap_thick_poly_0[3|2]/vout fgcell_amp_MOS_cap_thick_poly_0[3|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|2]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|2] fgcell_amp_MOS_cap_thick_poly_0[4|2]/vout fgcell_amp_MOS_cap_thick_poly_0[4|2]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|2]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|2]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|2]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|2]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|3] fgcell_amp_MOS_cap_thick_poly_0[0|3]/vout fgcell_amp_MOS_cap_thick_poly_0[0|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|3]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|3] fgcell_amp_MOS_cap_thick_poly_0[1|3]/vout fgcell_amp_MOS_cap_thick_poly_0[1|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|3]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|3] fgcell_amp_MOS_cap_thick_poly_0[2|3]/vout fgcell_amp_MOS_cap_thick_poly_0[2|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|3]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|3] fgcell_amp_MOS_cap_thick_poly_0[3|3]/vout fgcell_amp_MOS_cap_thick_poly_0[3|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|3]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|3] fgcell_amp_MOS_cap_thick_poly_0[4|3]/vout fgcell_amp_MOS_cap_thick_poly_0[4|3]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|3]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|3]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|3]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|3]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|4] fgcell_amp_MOS_cap_thick_poly_0[0|4]/vout fgcell_amp_MOS_cap_thick_poly_0[0|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|4]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|4]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|4] fgcell_amp_MOS_cap_thick_poly_0[1|4]/vout fgcell_amp_MOS_cap_thick_poly_0[1|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|4]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|4]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|4] fgcell_amp_MOS_cap_thick_poly_0[2|4]/vout fgcell_amp_MOS_cap_thick_poly_0[2|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|4]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|4]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|4] fgcell_amp_MOS_cap_thick_poly_0[3|4]/vout fgcell_amp_MOS_cap_thick_poly_0[3|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|4]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|4]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|4] fgcell_amp_MOS_cap_thick_poly_0[4|4]/vout fgcell_amp_MOS_cap_thick_poly_0[4|4]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|4]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|4]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|4]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|4]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|5] fgcell_amp_MOS_cap_thick_poly_0[0|5]/vout fgcell_amp_MOS_cap_thick_poly_0[0|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|5]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|5] fgcell_amp_MOS_cap_thick_poly_0[1|5]/vout fgcell_amp_MOS_cap_thick_poly_0[1|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|5]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|5] fgcell_amp_MOS_cap_thick_poly_0[2|5]/vout fgcell_amp_MOS_cap_thick_poly_0[2|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|5]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|5] fgcell_amp_MOS_cap_thick_poly_0[3|5]/vout fgcell_amp_MOS_cap_thick_poly_0[3|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|5]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|5] fgcell_amp_MOS_cap_thick_poly_0[4|5]/vout fgcell_amp_MOS_cap_thick_poly_0[4|5]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|5]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|5]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|5]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|5]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|6] fgcell_amp_MOS_cap_thick_poly_0[0|6]/vout fgcell_amp_MOS_cap_thick_poly_0[0|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|6]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|6] fgcell_amp_MOS_cap_thick_poly_0[1|6]/vout fgcell_amp_MOS_cap_thick_poly_0[1|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|6]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|6] fgcell_amp_MOS_cap_thick_poly_0[2|6]/vout fgcell_amp_MOS_cap_thick_poly_0[2|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|6]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|6] fgcell_amp_MOS_cap_thick_poly_0[3|6]/vout fgcell_amp_MOS_cap_thick_poly_0[3|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|6]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|6] fgcell_amp_MOS_cap_thick_poly_0[4|6]/vout fgcell_amp_MOS_cap_thick_poly_0[4|6]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|6]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|6]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|6]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|6]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|7] fgcell_amp_MOS_cap_thick_poly_0[0|7]/vout fgcell_amp_MOS_cap_thick_poly_0[0|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|7]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|7] fgcell_amp_MOS_cap_thick_poly_0[1|7]/vout fgcell_amp_MOS_cap_thick_poly_0[1|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|7]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|7] fgcell_amp_MOS_cap_thick_poly_0[2|7]/vout fgcell_amp_MOS_cap_thick_poly_0[2|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|7]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|7] fgcell_amp_MOS_cap_thick_poly_0[3|7]/vout fgcell_amp_MOS_cap_thick_poly_0[3|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|7]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|7] fgcell_amp_MOS_cap_thick_poly_0[4|7]/vout fgcell_amp_MOS_cap_thick_poly_0[4|7]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|7]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|7]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|7]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|7]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|8] fgcell_amp_MOS_cap_thick_poly_0[0|8]/vout fgcell_amp_MOS_cap_thick_poly_0[0|8]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|8]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|8] fgcell_amp_MOS_cap_thick_poly_0[1|8]/vout fgcell_amp_MOS_cap_thick_poly_0[1|8]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|8]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|8] fgcell_amp_MOS_cap_thick_poly_0[2|8]/vout fgcell_amp_MOS_cap_thick_poly_0[2|8]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|8]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|8] fgcell_amp_MOS_cap_thick_poly_0[3|8]/vout fgcell_amp_MOS_cap_thick_poly_0[3|8]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|8]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|8] fgcell_amp_MOS_cap_thick_poly_0[4|8]/vout fgcell_amp_MOS_cap_thick_poly_0[4|8]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|8]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|8]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|8]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|8]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[0|9] fgcell_amp_MOS_cap_thick_poly_0[0|9]/vout fgcell_amp_MOS_cap_thick_poly_0[0|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[0|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[0|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[0|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[0|9]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[1|9] fgcell_amp_MOS_cap_thick_poly_0[1|9]/vout fgcell_amp_MOS_cap_thick_poly_0[1|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[1|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[1|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[1|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[1|9]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[2|9] fgcell_amp_MOS_cap_thick_poly_0[2|9]/vout fgcell_amp_MOS_cap_thick_poly_0[2|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[2|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[2|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[2|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[2|9]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[3|9] fgcell_amp_MOS_cap_thick_poly_0[3|9]/vout fgcell_amp_MOS_cap_thick_poly_0[3|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[3|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[3|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[3|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[3|9]/vinj fgcell_amp_MOS_cap_thick_poly
Xfgcell_amp_MOS_cap_thick_poly_0[4|9] fgcell_amp_MOS_cap_thick_poly_0[4|9]/vout fgcell_amp_MOS_cap_thick_poly_0[4|9]/vdd
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/row_en_b fgcell_amp_MOS_cap_thick_poly_0[4|9]/x1/vtun
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/VSRC fgcell_amp_MOS_cap_thick_poly_0[4|9]/x1/vctrl
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/row_en VSUBS fgcell_amp_MOS_cap_thick_poly_0[4|9]/x2/vb
+ fgcell_amp_MOS_cap_thick_poly_0[4|9]/vinj fgcell_amp_MOS_cap_thick_poly
.ends

.subckt array_row_decode a[4] a[3] a[2] a[1] a[0] w[31] w[30] w[29] w[28] w[27] w[26]
+ w[25] w[24] w[23] w[22] w[21] w[20] w[19] w[18] w[17] w[16] w[15] w[14] w[13] w[12]
+ w[11] w[10] w[9] w[8] w[7] w[6] w[5] w[4] w[3] w[2] w[1] w[0] VGND VPWR
Xx1 a[4] VGND VGND VPWR VPWR x1/Y sky130_fd_sc_hd__inv_1
Xx3 a[2] VGND VGND VPWR VPWR x3/Y sky130_fd_sc_hd__inv_1
Xx2 a[3] VGND VGND VPWR VPWR x2/Y sky130_fd_sc_hd__inv_1
Xx4 a[1] VGND VGND VPWR VPWR x6/B sky130_fd_sc_hd__inv_1
Xx5 a[0] VGND VGND VPWR VPWR x8/A sky130_fd_sc_hd__inv_1
Xx6 x8/A x6/B VGND VGND VPWR VPWR x6/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand2_2_0 a[0] x6/B VGND VGND VPWR VPWR sky130_fd_sc_hd__nand2_2_0/Y
+ sky130_fd_sc_hd__nand2_2
Xx8 x8/A a[1] VGND VGND VPWR VPWR x8/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_1[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xx9 a[0] a[1] VGND VGND VPWR VPWR x9/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__decap_3_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xx10 x3/Y x2/Y VGND VGND VPWR VPWR x10/Y sky130_fd_sc_hd__nand2_2
Xx11 a[2] x2/Y VGND VGND VPWR VPWR x11/Y sky130_fd_sc_hd__nand2_2
Xx12 x3/Y a[3] VGND VGND VPWR VPWR x12/Y sky130_fd_sc_hd__nand2_2
Xx13 a[2] a[3] VGND VGND VPWR VPWR x13/Y sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nor3_1_0[0] x8/Y x13/Y x1/Y VGND VGND VPWR VPWR w[30] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[1] x6/Y x13/Y x1/Y VGND VGND VPWR VPWR w[28] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[2] x8/Y x12/Y x1/Y VGND VGND VPWR VPWR w[26] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[3] x6/Y x12/Y x1/Y VGND VGND VPWR VPWR w[24] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[4] x8/Y x11/Y x1/Y VGND VGND VPWR VPWR w[22] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[5] x6/Y x11/Y x1/Y VGND VGND VPWR VPWR w[20] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[6] x8/Y x10/Y x1/Y VGND VGND VPWR VPWR w[18] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[7] x6/Y x10/Y x1/Y VGND VGND VPWR VPWR w[16] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[8] x8/Y x13/Y a[4] VGND VGND VPWR VPWR w[14] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[9] x6/Y x13/Y a[4] VGND VGND VPWR VPWR w[12] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[10] x8/Y x12/Y a[4] VGND VGND VPWR VPWR w[10] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[11] x6/Y x12/Y a[4] VGND VGND VPWR VPWR w[8] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[12] x8/Y x11/Y a[4] VGND VGND VPWR VPWR w[6] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[13] x6/Y x11/Y a[4] VGND VGND VPWR VPWR w[4] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[14] x8/Y x10/Y a[4] VGND VGND VPWR VPWR w[2] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_0[15] x6/Y x10/Y a[4] VGND VGND VPWR VPWR w[0] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[0] x9/Y x13/Y x1/Y VGND VGND VPWR VPWR w[31] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[1] sky130_fd_sc_hd__nand2_2_0/Y x13/Y x1/Y VGND VGND VPWR
+ VPWR w[29] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[2] x9/Y x12/Y x1/Y VGND VGND VPWR VPWR w[27] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[3] sky130_fd_sc_hd__nand2_2_0/Y x12/Y x1/Y VGND VGND VPWR
+ VPWR w[25] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[4] x9/Y x11/Y x1/Y VGND VGND VPWR VPWR w[23] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[5] sky130_fd_sc_hd__nand2_2_0/Y x11/Y x1/Y VGND VGND VPWR
+ VPWR w[21] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[6] x9/Y x10/Y x1/Y VGND VGND VPWR VPWR w[19] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[7] sky130_fd_sc_hd__nand2_2_0/Y x10/Y x1/Y VGND VGND VPWR
+ VPWR w[17] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[8] x9/Y x13/Y a[4] VGND VGND VPWR VPWR w[15] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[9] sky130_fd_sc_hd__nand2_2_0/Y x13/Y a[4] VGND VGND VPWR
+ VPWR w[13] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[10] x9/Y x12/Y a[4] VGND VGND VPWR VPWR w[11] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[11] sky130_fd_sc_hd__nand2_2_0/Y x12/Y a[4] VGND VGND VPWR
+ VPWR w[9] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[12] x9/Y x11/Y a[4] VGND VGND VPWR VPWR w[7] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[13] sky130_fd_sc_hd__nand2_2_0/Y x11/Y a[4] VGND VGND VPWR
+ VPWR w[5] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[14] x9/Y x10/Y a[4] VGND VGND VPWR VPWR w[3] sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_1_1[15] sky130_fd_sc_hd__nand2_2_0/Y x10/Y a[4] VGND VGND VPWR
+ VPWR w[1] sky130_fd_sc_hd__nor3_1
.ends

.subckt fgcell_amp x1/vtun tg5v0_0/vout x2/VDD x2/v1 x1/vinj_en_b x1/vsrc x1/vctrl
+ tg5v0_0/en VSUBS x1/vinj x2/vb
Xx1 x1/vinj x1/vinj_en_b x1/vtun x1/vctrl x1/vsrc VSUBS x2/v1 fgcell
Xx2 x2/v1 x2/v2 VSUBS x2/VDD x2/vb x2/v2 diffamp_nmos
Xtg5v0_0 x2/v2 tg5v0_0/vout tg5v0_0/en x1/vinj_en_b x1/vinj VSUBS tg5v0
.ends

.subckt fgcell_amp_MiM_cap_1_5 vinj vtun x1/tg5v0_0/vout row_en x1/x1/vctrl x1/x2/vb
+ vdd vsrc row_en_b VGND
Xx1 vtun x1/tg5v0_0/vout vdd x1/x2/v1 row_en vsrc x1/x1/vctrl row_en_b VGND vinj x1/x2/vb
+ fgcell_amp
X0 x1/x2/v1 VGND sky130_fd_pr__cap_mim_m3_1 l=1 w=5
.ends

.subckt array_core_block1 fgcell_amp_MiM_cap_1_5_0[7|7]/vtun fgcell_amp_MiM_cap_1_5_0[0|3]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[8|5]/vsrc fgcell_amp_MiM_cap_1_5_0[9|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[5|9]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[6|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[5|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|4]/vinj
+ fgcell_amp_MiM_cap_1_5_0[9|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|9]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|4]/vsrc fgcell_amp_MiM_cap_1_5_0[2|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[3|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|5]/vinj fgcell_amp_MiM_cap_1_5_0[2|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|0]/vsrc fgcell_amp_MiM_cap_1_5_0[0|5]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[8|7]/vsrc fgcell_amp_MiM_cap_1_5_0[6|6]/vdd fgcell_amp_MiM_cap_1_5_0[4|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|3]/vtun fgcell_amp_MiM_cap_1_5_0[2|6]/vinj fgcell_amp_MiM_cap_1_5_0[3|1]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[8|6]/vsrc fgcell_amp_MiM_cap_1_5_0[9|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[0|6]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[8|8]/vsrc fgcell_amp_MiM_cap_1_5_0[5|4]/vdd fgcell_amp_MiM_cap_1_5_0[6|7]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[5|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[9|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|1]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[5|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|7]/vinj
+ fgcell_amp_MiM_cap_1_5_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|4]/vtun fgcell_amp_MiM_cap_1_5_0[3|2]/vsrc fgcell_amp_MiM_cap_1_5_0[0|4]/vdd
+ fgcell_amp_MiM_cap_1_5_0[0|7]/vsrc fgcell_amp_MiM_cap_1_5_0[2|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|9]/vsrc fgcell_amp_MiM_cap_1_5_0[8|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|8]/vinj fgcell_amp_MiM_cap_1_5_0[5|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|3]/vsrc fgcell_amp_MiM_cap_1_5_0[0|8]/vsrc fgcell_amp_MiM_cap_1_5_0[4|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[9|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|4]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[0|9]/vsrc fgcell_amp_MiM_cap_1_5_0[7|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|0]/vinj fgcell_amp_MiM_cap_1_5_0[0|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|2]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[7|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|7]/vtun fgcell_amp_MiM_cap_1_5_0[6|0]/vsrc fgcell_amp_MiM_cap_1_5_0[4|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|5]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[1|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|5]/vsrc fgcell_amp_MiM_cap_1_5_0[0|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[5|5]/vdd fgcell_amp_MiM_cap_1_5_0[8|1]/vinj
+ fgcell_amp_MiM_cap_1_5_0[3|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|3]/vdd
+ fgcell_amp_MiM_cap_1_5_0[9|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|1]/vsrc fgcell_amp_MiM_cap_1_5_0[8|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|0]/vinj
+ fgcell_amp_MiM_cap_1_5_0[8|2]/vinj fgcell_amp_MiM_cap_1_5_0[2|9]/vdd fgcell_amp_MiM_cap_1_5_0[9|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|2]/vsrc fgcell_amp_MiM_cap_1_5_0[3|7]/vsrc fgcell_amp_MiM_cap_1_5_0[7|9]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[6|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|1]/vinj fgcell_amp_MiM_cap_1_5_0[5|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|3]/vinj fgcell_amp_MiM_cap_1_5_0[2|9]/row_en_b fgcell_amp_MiM_cap_1_5_0[6|0]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[2|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|3]/vsrc fgcell_amp_MiM_cap_1_5_0[3|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|8]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[0|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|2]/vinj fgcell_amp_MiM_cap_1_5_0[6|8]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[5|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|4]/vinj fgcell_amp_MiM_cap_1_5_0[8|1]/vtun fgcell_amp_MiM_cap_1_5_0[3|0]/vdd
+ fgcell_amp_MiM_cap_1_5_0[0|3]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[9|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|9]/vtun fgcell_amp_MiM_cap_1_5_0[6|4]/vsrc fgcell_amp_MiM_cap_1_5_0[3|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|8]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|3]/vinj fgcell_amp_MiM_cap_1_5_0[5|6]/vdd
+ fgcell_amp_MiM_cap_1_5_0[8|5]/vinj fgcell_amp_MiM_cap_1_5_0[5|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|0]/vtun fgcell_amp_MiM_cap_1_5_0[8|2]/vtun fgcell_amp_MiM_cap_1_5_0[9|0]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[1|3]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[6|5]/vsrc fgcell_amp_MiM_cap_1_5_0[5|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|4]/vinj
+ fgcell_amp_MiM_cap_1_5_0[6|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[0|1]/vtun fgcell_amp_MiM_cap_1_5_0[8|6]/vinj fgcell_amp_MiM_cap_1_5_0[8|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[8|3]/vtun fgcell_amp_MiM_cap_1_5_0[3|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|1]/vsrc fgcell_amp_MiM_cap_1_5_0[1|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|4]/vdd fgcell_amp_MiM_cap_1_5_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|0]/vinj fgcell_amp_MiM_cap_1_5_0[8|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|5]/vinj fgcell_amp_MiM_cap_1_5_0[8|7]/vinj
+ fgcell_amp_MiM_cap_1_5_0[7|9]/vdd fgcell_amp_MiM_cap_1_5_0[0|2]/vtun fgcell_amp_MiM_cap_1_5_0[8|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|0]/vsrc fgcell_amp_MiM_cap_1_5_0[9|2]/vsrc fgcell_amp_MiM_cap_1_5_0[3|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|7]/vsrc fgcell_amp_MiM_cap_1_5_0[4|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|5]/vdd fgcell_amp_MiM_cap_1_5_0[3|1]/vinj
+ fgcell_amp_MiM_cap_1_5_0[5|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|6]/vinj fgcell_amp_MiM_cap_1_5_0[4|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|3]/vtun fgcell_amp_MiM_cap_1_5_0[6|9]/vdd fgcell_amp_MiM_cap_1_5_0[8|8]/vinj
+ fgcell_amp_MiM_cap_1_5_0[8|5]/vtun fgcell_amp_MiM_cap_1_5_0[1|1]/vsrc fgcell_amp_MiM_cap_1_5_0[4|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|3]/vsrc fgcell_amp_MiM_cap_1_5_0[6|8]/vsrc fgcell_amp_MiM_cap_1_5_0[9|5]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[5|0]/vinj fgcell_amp_MiM_cap_1_5_0[6|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|7]/vinj fgcell_amp_MiM_cap_1_5_0[5|7]/vdd
+ fgcell_amp_MiM_cap_1_5_0[8|0]/vdd fgcell_amp_MiM_cap_1_5_0[0|4]/vtun fgcell_amp_MiM_cap_1_5_0[4|5]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[1|2]/vsrc fgcell_amp_MiM_cap_1_5_0[9|4]/vsrc fgcell_amp_MiM_cap_1_5_0[5|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|0]/vtun fgcell_amp_MiM_cap_1_5_0[0|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|8]/vinj fgcell_amp_MiM_cap_1_5_0[4|1]/vdd
+ fgcell_amp_MiM_cap_1_5_0[0|5]/vtun fgcell_amp_MiM_cap_1_5_0[8|7]/vtun fgcell_amp_MiM_cap_1_5_0[1|3]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[1|9]/vdd fgcell_amp_MiM_cap_1_5_0[8|3]/vdd fgcell_amp_MiM_cap_1_5_0[6|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|5]/vsrc fgcell_amp_MiM_cap_1_5_0[5|1]/vinj fgcell_amp_MiM_cap_1_5_0[3|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[1|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|4]/vinj fgcell_amp_MiM_cap_1_5_0[3|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|6]/vtun fgcell_amp_MiM_cap_1_5_0[3|3]/vdd fgcell_amp_MiM_cap_1_5_0[3|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[8|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|9]/vinj fgcell_amp_MiM_cap_1_5_0[0|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|8]/vtun fgcell_amp_MiM_cap_1_5_0[1|4]/vsrc fgcell_amp_MiM_cap_1_5_0[9|6]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[7|3]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[6|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|9]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|4]/vdd fgcell_amp_MiM_cap_1_5_0[7|6]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[5|0]/vtun fgcell_amp_MiM_cap_1_5_0[3|5]/vinj fgcell_amp_MiM_cap_1_5_0[5|2]/vinj
+ fgcell_amp_MiM_cap_1_5_0[6|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|9]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[9|7]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|0]/vsrc fgcell_amp_MiM_cap_1_5_0[1|3]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[0|7]/vtun fgcell_amp_MiM_cap_1_5_0[5|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|5]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|0]/vdd fgcell_amp_MiM_cap_1_5_0[8|3]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[9|7]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[5|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|0]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[8|9]/vinj fgcell_amp_MiM_cap_1_5_0[2|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|6]/vinj fgcell_amp_MiM_cap_1_5_0[3|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|1]/vsrc fgcell_amp_MiM_cap_1_5_0[2|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|8]/vdd fgcell_amp_MiM_cap_1_5_0[1|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|6]/vsrc fgcell_amp_MiM_cap_1_5_0[9|8]/vsrc fgcell_amp_MiM_cap_1_5_0[9|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|6]/vdd fgcell_amp_MiM_cap_1_5_0[2|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[5|1]/vtun fgcell_amp_MiM_cap_1_5_0[8|4]/row_en fgcell_amp_MiM_cap_1_5_0[1|6]/vdd
+ fgcell_amp_MiM_cap_1_5_0[5|3]/vinj fgcell_amp_MiM_cap_1_5_0[5|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|4]/row_en fgcell_amp_MiM_cap_1_5_0[0|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|7]/vinj
+ fgcell_amp_MiM_cap_1_5_0[3|4]/vtun fgcell_amp_MiM_cap_1_5_0[0|8]/vdd fgcell_amp_MiM_cap_1_5_0[4|2]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[0|9]/vtun fgcell_amp_MiM_cap_1_5_0[1|7]/vsrc fgcell_amp_MiM_cap_1_5_0[9|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[5|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|5]/row_en fgcell_amp_MiM_cap_1_5_0[1|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|8]/vinj
+ fgcell_amp_MiM_cap_1_5_0[5|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|5]/vtun fgcell_amp_MiM_cap_1_5_0[5|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|3]/vsrc fgcell_amp_MiM_cap_1_5_0[3|4]/vdd fgcell_amp_MiM_cap_1_5_0[5|4]/vinj
+ fgcell_amp_MiM_cap_1_5_0[6|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[0|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[9|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|8]/vsrc fgcell_amp_MiM_cap_1_5_0[7|2]/vdd fgcell_amp_MiM_cap_1_5_0[3|4]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[4|0]/row_en fgcell_amp_MiM_cap_1_5_0[8|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|1]/vtun fgcell_amp_MiM_cap_1_5_0[8|9]/vtun fgcell_amp_MiM_cap_1_5_0[7|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|9]/vinj fgcell_amp_MiM_cap_1_5_0[0|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[9|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|6]/vtun fgcell_amp_MiM_cap_1_5_0[8|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|4]/vsrc fgcell_amp_MiM_cap_1_5_0[2|2]/vdd fgcell_amp_MiM_cap_1_5_0[1|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|6]/row_en fgcell_amp_MiM_cap_1_5_0[1|9]/vsrc fgcell_amp_MiM_cap_1_5_0[1|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|1]/row_en fgcell_amp_MiM_cap_1_5_0[5|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|0]/vinj fgcell_amp_MiM_cap_1_5_0[5|5]/vinj fgcell_amp_MiM_cap_1_5_0[4|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|1]/row_en fgcell_amp_MiM_cap_1_5_0[3|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|0]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[3|7]/vtun fgcell_amp_MiM_cap_1_5_0[7|0]/vdd fgcell_amp_MiM_cap_1_5_0[4|5]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|4]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|9]/vdd fgcell_amp_MiM_cap_1_5_0[3|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|7]/vdd fgcell_amp_MiM_cap_1_5_0[9|1]/vinj fgcell_amp_MiM_cap_1_5_0[7|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|2]/row_en fgcell_amp_MiM_cap_1_5_0[6|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|1]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[6|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|8]/vtun fgcell_amp_MiM_cap_1_5_0[3|1]/vdd
+ fgcell_amp_MiM_cap_1_5_0[4|6]/vsrc fgcell_amp_MiM_cap_1_5_0[0|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[3|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[3|4]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|9]/vdd fgcell_amp_MiM_cap_1_5_0[4|7]/vdd fgcell_amp_MiM_cap_1_5_0[6|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|6]/vinj fgcell_amp_MiM_cap_1_5_0[7|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[6|6]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[1|0]/vinj fgcell_amp_MiM_cap_1_5_0[9|2]/vinj fgcell_amp_MiM_cap_1_5_0[2|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|3]/row_en fgcell_amp_MiM_cap_1_5_0[6|4]/vtun fgcell_amp_MiM_cap_1_5_0[5|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|2]/vsrc fgcell_amp_MiM_cap_1_5_0[3|9]/vtun fgcell_amp_MiM_cap_1_5_0[3|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[5|9]/row_en fgcell_amp_MiM_cap_1_5_0[8|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|7]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[4|4]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[9|9]/row_en fgcell_amp_MiM_cap_1_5_0[7|3]/vdd
+ fgcell_amp_MiM_cap_1_5_0[3|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[1|1]/vinj fgcell_amp_MiM_cap_1_5_0[9|3]/vinj fgcell_amp_MiM_cap_1_5_0[8|4]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|9]/row_en fgcell_amp_MiM_cap_1_5_0[9|0]/vtun fgcell_amp_MiM_cap_1_5_0[5|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|5]/vtun fgcell_amp_MiM_cap_1_5_0[9|4]/row_en fgcell_amp_MiM_cap_1_5_0[6|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|3]/vsrc fgcell_amp_MiM_cap_1_5_0[5|7]/vinj fgcell_amp_MiM_cap_1_5_0[4|8]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[2|3]/vdd fgcell_amp_MiM_cap_1_5_0[6|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[5|4]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|0]/vdd fgcell_amp_MiM_cap_1_5_0[6|0]/vinj
+ fgcell_amp_MiM_cap_1_5_0[2|4]/row_en fgcell_amp_MiM_cap_1_5_0[6|1]/vdd fgcell_amp_MiM_cap_1_5_0[4|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|2]/vinj fgcell_amp_MiM_cap_1_5_0[4|5]/vdd
+ fgcell_amp_MiM_cap_1_5_0[9|4]/vinj fgcell_amp_MiM_cap_1_5_0[6|9]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|5]/row_en fgcell_amp_MiM_cap_1_5_0[9|1]/vtun fgcell_amp_MiM_cap_1_5_0[6|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|8]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|4]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[1|5]/row_en fgcell_amp_MiM_cap_1_5_0[4|6]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[5|5]/row_en fgcell_amp_MiM_cap_1_5_0[6|4]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[8|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[5|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|6]/vdd fgcell_amp_MiM_cap_1_5_0[5|8]/vinj
+ fgcell_amp_MiM_cap_1_5_0[2|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[5|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|3]/vinj fgcell_amp_MiM_cap_1_5_0[9|5]/vinj
+ fgcell_amp_MiM_cap_1_5_0[1|0]/vtun fgcell_amp_MiM_cap_1_5_0[9|2]/vtun fgcell_amp_MiM_cap_1_5_0[1|8]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[6|1]/vinj fgcell_amp_MiM_cap_1_5_0[5|0]/row_en fgcell_amp_MiM_cap_1_5_0[9|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|7]/vtun fgcell_amp_MiM_cap_1_5_0[0|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|5]/vsrc fgcell_amp_MiM_cap_1_5_0[9|8]/vdd fgcell_amp_MiM_cap_1_5_0[4|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|6]/row_en fgcell_amp_MiM_cap_1_5_0[4|8]/vdd fgcell_amp_MiM_cap_1_5_0[2|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[5|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[8|6]/vdd fgcell_amp_MiM_cap_1_5_0[1|4]/vinj
+ fgcell_amp_MiM_cap_1_5_0[1|6]/row_en fgcell_amp_MiM_cap_1_5_0[1|1]/vtun fgcell_amp_MiM_cap_1_5_0[9|6]/vinj
+ fgcell_amp_MiM_cap_1_5_0[4|1]/row_en fgcell_amp_MiM_cap_1_5_0[2|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|3]/vtun fgcell_amp_MiM_cap_1_5_0[8|1]/row_en fgcell_amp_MiM_cap_1_5_0[6|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|1]/vdd fgcell_amp_MiM_cap_1_5_0[1|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|7]/vtun fgcell_amp_MiM_cap_1_5_0[7|7]/row_en fgcell_amp_MiM_cap_1_5_0[5|9]/vinj
+ fgcell_amp_MiM_cap_1_5_0[5|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|6]/vdd fgcell_amp_MiM_cap_1_5_0[0|7]/row_en fgcell_amp_MiM_cap_1_5_0[7|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|0]/vinj fgcell_amp_MiM_cap_1_5_0[6|2]/vinj fgcell_amp_MiM_cap_1_5_0[4|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|5]/vinj fgcell_amp_MiM_cap_1_5_0[9|7]/vinj fgcell_amp_MiM_cap_1_5_0[7|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|2]/vtun fgcell_amp_MiM_cap_1_5_0[9|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|0]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[4|2]/vdd fgcell_amp_MiM_cap_1_5_0[8|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|7]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[0|2]/row_en fgcell_amp_MiM_cap_1_5_0[5|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|4]/vdd fgcell_amp_MiM_cap_1_5_0[2|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|0]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[3|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[9|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[6|2]/vdd fgcell_amp_MiM_cap_1_5_0[1|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[3|8]/row_en fgcell_amp_MiM_cap_1_5_0[8|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|1]/vinj
+ fgcell_amp_MiM_cap_1_5_0[1|0]/row_en fgcell_amp_MiM_cap_1_5_0[3|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[5|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|6]/vinj fgcell_amp_MiM_cap_1_5_0[7|8]/row_en fgcell_amp_MiM_cap_1_5_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|8]/vinj fgcell_amp_MiM_cap_1_5_0[0|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|1]/vsrc fgcell_amp_MiM_cap_1_5_0[0|3]/vdd fgcell_amp_MiM_cap_1_5_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|8]/vsrc fgcell_amp_MiM_cap_1_5_0[6|0]/vdd fgcell_amp_MiM_cap_1_5_0[6|3]/vinj
+ fgcell_amp_MiM_cap_1_5_0[1|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[9|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[1|2]/vdd fgcell_amp_MiM_cap_1_5_0[7|3]/row_en fgcell_amp_MiM_cap_1_5_0[9|5]/vdd
+ fgcell_amp_MiM_cap_1_5_0[6|9]/row_en fgcell_amp_MiM_cap_1_5_0[9|0]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|2]/vinj fgcell_amp_MiM_cap_1_5_0[4|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|3]/row_en fgcell_amp_MiM_cap_1_5_0[1|7]/vinj fgcell_amp_MiM_cap_1_5_0[9|9]/vinj
+ fgcell_amp_MiM_cap_1_5_0[1|4]/vtun fgcell_amp_MiM_cap_1_5_0[9|6]/vtun fgcell_amp_MiM_cap_1_5_0[1|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|2]/vsrc fgcell_amp_MiM_cap_1_5_0[3|9]/row_en fgcell_amp_MiM_cap_1_5_0[7|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[6|4]/row_en fgcell_amp_MiM_cap_1_5_0[0|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|1]/vdd
+ fgcell_amp_MiM_cap_1_5_0[4|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|3]/vinj fgcell_amp_MiM_cap_1_5_0[4|0]/vtun fgcell_amp_MiM_cap_1_5_0[6|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|8]/vinj fgcell_amp_MiM_cap_1_5_0[6|4]/vinj fgcell_amp_MiM_cap_1_5_0[8|7]/vdd
+ fgcell_amp_MiM_cap_1_5_0[8|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|5]/vtun fgcell_amp_MiM_cap_1_5_0[9|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|3]/vsrc fgcell_amp_MiM_cap_1_5_0[0|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|9]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[4|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[1|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[3|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[0|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|7]/vdd
+ fgcell_amp_MiM_cap_1_5_0[1|7]/vdd fgcell_amp_MiM_cap_1_5_0[2|5]/row_en fgcell_amp_MiM_cap_1_5_0[0|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|4]/vinj fgcell_amp_MiM_cap_1_5_0[0|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|5]/vdd fgcell_amp_MiM_cap_1_5_0[7|4]/vdd fgcell_amp_MiM_cap_1_5_0[6|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|9]/vinj fgcell_amp_MiM_cap_1_5_0[1|2]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|6]/vtun fgcell_amp_MiM_cap_1_5_0[9|8]/vtun fgcell_amp_MiM_cap_1_5_0[3|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|4]/vsrc fgcell_amp_MiM_cap_1_5_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|0]/row_en fgcell_amp_MiM_cap_1_5_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|0]/vdd fgcell_amp_MiM_cap_1_5_0[6|5]/vinj fgcell_amp_MiM_cap_1_5_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|6]/row_en fgcell_amp_MiM_cap_1_5_0[4|5]/vinj
+ fgcell_amp_MiM_cap_1_5_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|5]/vdd fgcell_amp_MiM_cap_1_5_0[6|3]/vdd fgcell_amp_MiM_cap_1_5_0[9|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|7]/vtun fgcell_amp_MiM_cap_1_5_0[5|0]/vsrc fgcell_amp_MiM_cap_1_5_0[9|2]/vdd
+ fgcell_amp_MiM_cap_1_5_0[8|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[9|9]/vtun fgcell_amp_MiM_cap_1_5_0[2|5]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[4|9]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|6]/vsrc fgcell_amp_MiM_cap_1_5_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|1]/row_en fgcell_amp_MiM_cap_1_5_0[3|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|1]/row_en fgcell_amp_MiM_cap_1_5_0[2|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|3]/vdd
+ fgcell_amp_MiM_cap_1_5_0[8|9]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|7]/row_en fgcell_amp_MiM_cap_1_5_0[4|6]/vinj
+ fgcell_amp_MiM_cap_1_5_0[5|1]/vdd fgcell_amp_MiM_cap_1_5_0[2|1]/row_en fgcell_amp_MiM_cap_1_5_0[6|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|3]/vtun fgcell_amp_MiM_cap_1_5_0[5|1]/vsrc fgcell_amp_MiM_cap_1_5_0[9|3]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[1|8]/vtun fgcell_amp_MiM_cap_1_5_0[1|7]/row_en fgcell_amp_MiM_cap_1_5_0[5|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|6]/vsrc fgcell_amp_MiM_cap_1_5_0[6|6]/vinj fgcell_amp_MiM_cap_1_5_0[6|6]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[5|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|6]/vsrc fgcell_amp_MiM_cap_1_5_0[5|7]/row_en fgcell_amp_MiM_cap_1_5_0[8|4]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[6|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|9]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[7|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|2]/row_en fgcell_amp_MiM_cap_1_5_0[4|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|3]/row_en_b fgcell_amp_MiM_cap_1_5_0[0|1]/vdd fgcell_amp_MiM_cap_1_5_0[3|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|2]/row_en fgcell_amp_MiM_cap_1_5_0[4|7]/vinj fgcell_amp_MiM_cap_1_5_0[1|6]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[9|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|2]/row_en fgcell_amp_MiM_cap_1_5_0[8|8]/vdd fgcell_amp_MiM_cap_1_5_0[2|0]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|9]/vtun fgcell_amp_MiM_cap_1_5_0[5|2]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[4|8]/row_en fgcell_amp_MiM_cap_1_5_0[2|7]/vsrc fgcell_amp_MiM_cap_1_5_0[2|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|9]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|1]/vdd fgcell_amp_MiM_cap_1_5_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[4|9]/vdd fgcell_amp_MiM_cap_1_5_0[9|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|8]/row_en fgcell_amp_MiM_cap_1_5_0[8|0]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|3]/row_en fgcell_amp_MiM_cap_1_5_0[7|0]/vtun fgcell_amp_MiM_cap_1_5_0[3|8]/vdd
+ fgcell_amp_MiM_cap_1_5_0[6|7]/vinj fgcell_amp_MiM_cap_1_5_0[2|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[2|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|8]/vinj fgcell_amp_MiM_cap_1_5_0[8|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|5]/vtun fgcell_amp_MiM_cap_1_5_0[7|6]/vdd fgcell_amp_MiM_cap_1_5_0[5|3]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[7|0]/vinj fgcell_amp_MiM_cap_1_5_0[7|9]/row_en fgcell_amp_MiM_cap_1_5_0[7|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|6]/vtun fgcell_amp_MiM_cap_1_5_0[2|8]/vsrc fgcell_amp_MiM_cap_1_5_0[3|2]/vdd
+ fgcell_amp_MiM_cap_1_5_0[5|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[0|9]/row_en fgcell_amp_MiM_cap_1_5_0[6|7]/vdd
+ fgcell_amp_MiM_cap_1_5_0[4|9]/row_en fgcell_amp_MiM_cap_1_5_0[5|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|6]/vdd fgcell_amp_MiM_cap_1_5_0[9|7]/row_en_b fgcell_amp_MiM_cap_1_5_0[7|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|9]/vinj fgcell_amp_MiM_cap_1_5_0[5|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[4|6]/vtun fgcell_amp_MiM_cap_1_5_0[6|4]/vdd fgcell_amp_MiM_cap_1_5_0[1|9]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|4]/vsrc fgcell_amp_MiM_cap_1_5_0[0|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|9]/vsrc fgcell_amp_MiM_cap_1_5_0[8|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|9]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[6|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|4]/row_en fgcell_amp_MiM_cap_1_5_0[6|8]/vinj fgcell_amp_MiM_cap_1_5_0[4|7]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[7|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[5|0]/vdd fgcell_amp_MiM_cap_1_5_0[2|8]/vdd
+ fgcell_amp_MiM_cap_1_5_0[1|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|1]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[7|1]/vinj fgcell_amp_MiM_cap_1_5_0[6|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|4]/vdd
+ fgcell_amp_MiM_cap_1_5_0[7|5]/vinj fgcell_amp_MiM_cap_1_5_0[6|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|5]/vdd fgcell_amp_MiM_cap_1_5_0[2|4]/row_en_b fgcell_amp_MiM_cap_1_5_0[8|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[0|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[8|0]/vsrc fgcell_amp_MiM_cap_1_5_0[2|9]/vinj fgcell_amp_MiM_cap_1_5_0[5|2]/vdd
+ fgcell_amp_MiM_cap_1_5_0[4|7]/vtun fgcell_amp_MiM_cap_1_5_0[5|5]/vsrc fgcell_amp_MiM_cap_1_5_0[9|0]/vdd
+ fgcell_amp_MiM_cap_1_5_0[3|5]/row_en fgcell_amp_MiM_cap_1_5_0[0|1]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|9]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|2]/vinj fgcell_amp_MiM_cap_1_5_0[7|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[1|1]/vdd fgcell_amp_MiM_cap_1_5_0[8|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|5]/row_en fgcell_amp_MiM_cap_1_5_0[0|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[3|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|2]/vdd fgcell_amp_MiM_cap_1_5_0[3|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|3]/vtun fgcell_amp_MiM_cap_1_5_0[4|6]/vdd
+ fgcell_amp_MiM_cap_1_5_0[7|6]/vinj fgcell_amp_MiM_cap_1_5_0[4|0]/vdd fgcell_amp_MiM_cap_1_5_0[7|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|8]/vtun fgcell_amp_MiM_cap_1_5_0[8|1]/vsrc fgcell_amp_MiM_cap_1_5_0[6|9]/vinj
+ fgcell_amp_MiM_cap_1_5_0[5|6]/vsrc fgcell_amp_MiM_cap_1_5_0[8|9]/vdd fgcell_amp_MiM_cap_1_5_0[6|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|0]/row_en fgcell_amp_MiM_cap_1_5_0[4|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[7|2]/vinj fgcell_amp_MiM_cap_1_5_0[9|5]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[1|1]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[2|0]/vinj fgcell_amp_MiM_cap_1_5_0[3|6]/row_en fgcell_amp_MiM_cap_1_5_0[8|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|7]/vdd fgcell_amp_MiM_cap_1_5_0[7|7]/vinj fgcell_amp_MiM_cap_1_5_0[6|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|3]/vinj fgcell_amp_MiM_cap_1_5_0[0|0]/vsrc fgcell_amp_MiM_cap_1_5_0[8|2]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[3|9]/vdd fgcell_amp_MiM_cap_1_5_0[7|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[4|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|7]/vsrc fgcell_amp_MiM_cap_1_5_0[7|7]/vdd fgcell_amp_MiM_cap_1_5_0[8|2]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[9|7]/row_en fgcell_amp_MiM_cap_1_5_0[7|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|9]/vdd fgcell_amp_MiM_cap_1_5_0[3|1]/row_en fgcell_amp_MiM_cap_1_5_0[1|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|5]/row_en_b fgcell_amp_MiM_cap_1_5_0[2|7]/row_en fgcell_amp_MiM_cap_1_5_0[2|1]/vinj
+ fgcell_amp_MiM_cap_1_5_0[2|8]/row_en_b fgcell_amp_MiM_cap_1_5_0[0|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[1|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|7]/row_en fgcell_amp_MiM_cap_1_5_0[7|8]/vinj
+ fgcell_amp_MiM_cap_1_5_0[9|1]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[7|5]/vtun fgcell_amp_MiM_cap_1_5_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|2]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[0|1]/vsrc fgcell_amp_MiM_cap_1_5_0[2|7]/vdd fgcell_amp_MiM_cap_1_5_0[7|3]/vinj
+ fgcell_amp_MiM_cap_1_5_0[8|3]/vsrc fgcell_amp_MiM_cap_1_5_0[2|5]/vdd fgcell_amp_MiM_cap_1_5_0[0|5]/row_en_b
+ fgcell_amp_MiM_cap_1_5_0[2|9]/vtun fgcell_amp_MiM_cap_1_5_0[5|8]/vsrc fgcell_amp_MiM_cap_1_5_0[6|5]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|2]/row_en fgcell_amp_MiM_cap_1_5_0[8|2]/vdd fgcell_amp_MiM_cap_1_5_0[0|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[6|2]/row_en fgcell_amp_MiM_cap_1_5_0[0|6]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[3|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_5_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|8]/row_en fgcell_amp_MiM_cap_1_5_0[2|2]/vinj
+ fgcell_amp_MiM_cap_1_5_0[3|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|9]/vinj fgcell_amp_MiM_cap_1_5_0[7|6]/vtun fgcell_amp_MiM_cap_1_5_0[1|5]/vdd
+ fgcell_amp_MiM_cap_1_5_0[0|2]/vsrc fgcell_amp_MiM_cap_1_5_0[8|4]/vsrc fgcell_amp_MiM_cap_1_5_0[5|3]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|8]/row_en fgcell_amp_MiM_cap_1_5_0[6|9]/vtun fgcell_amp_MiM_cap_1_5_0[5|9]/vsrc
+ fgcell_amp_MiM_cap_1_5_0[4|3]/vdd fgcell_amp_MiM_cap_1_5_0[5|3]/row_en fgcell_amp_MiM_cap_1_5_0[3|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[9|1]/vdd VSUBS fgcell_amp_MiM_cap_1_5_0[9|3]/row_en fgcell_amp_MiM_cap_1_5_0[1|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|2]/vtun fgcell_amp_MiM_cap_1_5_0[7|4]/vinj fgcell_amp_MiM_cap_1_5_0[7|8]/vdd
+ fgcell_amp_MiM_cap_1_5_0[2|3]/vinj fgcell_amp_MiM_cap_1_5_0[6|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_5_0[8|9]/row_en fgcell_amp_MiM_cap_1_5_0[0|2]/x1/x2/vb fgcell_amp_MiM_cap_1_5_0[2|0]/vtun
Xfgcell_amp_MiM_cap_1_5_0[0|0] fgcell_amp_MiM_cap_1_5_0[0|0]/vinj fgcell_amp_MiM_cap_1_5_0[0|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|0]/vdd fgcell_amp_MiM_cap_1_5_0[0|0]/vsrc fgcell_amp_MiM_cap_1_5_0[0|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|0] fgcell_amp_MiM_cap_1_5_0[1|0]/vinj fgcell_amp_MiM_cap_1_5_0[1|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|0]/vdd fgcell_amp_MiM_cap_1_5_0[1|0]/vsrc fgcell_amp_MiM_cap_1_5_0[1|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|0] fgcell_amp_MiM_cap_1_5_0[2|0]/vinj fgcell_amp_MiM_cap_1_5_0[2|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|0]/vdd fgcell_amp_MiM_cap_1_5_0[2|0]/vsrc fgcell_amp_MiM_cap_1_5_0[2|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|0] fgcell_amp_MiM_cap_1_5_0[3|0]/vinj fgcell_amp_MiM_cap_1_5_0[3|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|0]/vdd fgcell_amp_MiM_cap_1_5_0[3|0]/vsrc fgcell_amp_MiM_cap_1_5_0[3|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|0] fgcell_amp_MiM_cap_1_5_0[4|0]/vinj fgcell_amp_MiM_cap_1_5_0[4|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|0]/vdd fgcell_amp_MiM_cap_1_5_0[4|0]/vsrc fgcell_amp_MiM_cap_1_5_0[4|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|0] fgcell_amp_MiM_cap_1_5_0[5|0]/vinj fgcell_amp_MiM_cap_1_5_0[5|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|0]/vdd fgcell_amp_MiM_cap_1_5_0[5|0]/vsrc fgcell_amp_MiM_cap_1_5_0[5|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|0] fgcell_amp_MiM_cap_1_5_0[6|0]/vinj fgcell_amp_MiM_cap_1_5_0[6|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|0]/vdd fgcell_amp_MiM_cap_1_5_0[6|0]/vsrc fgcell_amp_MiM_cap_1_5_0[6|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|0] fgcell_amp_MiM_cap_1_5_0[7|0]/vinj fgcell_amp_MiM_cap_1_5_0[7|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|0]/vdd fgcell_amp_MiM_cap_1_5_0[7|0]/vsrc fgcell_amp_MiM_cap_1_5_0[7|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|0] fgcell_amp_MiM_cap_1_5_0[8|0]/vinj fgcell_amp_MiM_cap_1_5_0[8|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|0]/vdd fgcell_amp_MiM_cap_1_5_0[8|0]/vsrc fgcell_amp_MiM_cap_1_5_0[8|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|0] fgcell_amp_MiM_cap_1_5_0[9|0]/vinj fgcell_amp_MiM_cap_1_5_0[9|0]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|0]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|0]/vdd fgcell_amp_MiM_cap_1_5_0[9|0]/vsrc fgcell_amp_MiM_cap_1_5_0[9|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|1] fgcell_amp_MiM_cap_1_5_0[0|1]/vinj fgcell_amp_MiM_cap_1_5_0[0|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|1]/vdd fgcell_amp_MiM_cap_1_5_0[0|1]/vsrc fgcell_amp_MiM_cap_1_5_0[0|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|1] fgcell_amp_MiM_cap_1_5_0[1|1]/vinj fgcell_amp_MiM_cap_1_5_0[1|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|1]/vdd fgcell_amp_MiM_cap_1_5_0[1|1]/vsrc fgcell_amp_MiM_cap_1_5_0[1|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|1] fgcell_amp_MiM_cap_1_5_0[2|1]/vinj fgcell_amp_MiM_cap_1_5_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|1]/vdd fgcell_amp_MiM_cap_1_5_0[2|1]/vsrc fgcell_amp_MiM_cap_1_5_0[2|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|1] fgcell_amp_MiM_cap_1_5_0[3|1]/vinj fgcell_amp_MiM_cap_1_5_0[3|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|1]/vdd fgcell_amp_MiM_cap_1_5_0[3|1]/vsrc fgcell_amp_MiM_cap_1_5_0[3|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|1] fgcell_amp_MiM_cap_1_5_0[4|1]/vinj fgcell_amp_MiM_cap_1_5_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|1]/vdd fgcell_amp_MiM_cap_1_5_0[4|1]/vsrc fgcell_amp_MiM_cap_1_5_0[4|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|1] fgcell_amp_MiM_cap_1_5_0[5|1]/vinj fgcell_amp_MiM_cap_1_5_0[5|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|1]/vdd fgcell_amp_MiM_cap_1_5_0[5|1]/vsrc fgcell_amp_MiM_cap_1_5_0[5|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|1] fgcell_amp_MiM_cap_1_5_0[6|1]/vinj fgcell_amp_MiM_cap_1_5_0[6|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|1]/vdd fgcell_amp_MiM_cap_1_5_0[6|1]/vsrc fgcell_amp_MiM_cap_1_5_0[6|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|1] fgcell_amp_MiM_cap_1_5_0[7|1]/vinj fgcell_amp_MiM_cap_1_5_0[7|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|1]/vdd fgcell_amp_MiM_cap_1_5_0[7|1]/vsrc fgcell_amp_MiM_cap_1_5_0[7|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|1] fgcell_amp_MiM_cap_1_5_0[8|1]/vinj fgcell_amp_MiM_cap_1_5_0[8|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|1]/vdd fgcell_amp_MiM_cap_1_5_0[8|1]/vsrc fgcell_amp_MiM_cap_1_5_0[8|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|1] fgcell_amp_MiM_cap_1_5_0[9|1]/vinj fgcell_amp_MiM_cap_1_5_0[9|1]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|1]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|1]/vdd fgcell_amp_MiM_cap_1_5_0[9|1]/vsrc fgcell_amp_MiM_cap_1_5_0[9|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|2] fgcell_amp_MiM_cap_1_5_0[0|2]/vinj fgcell_amp_MiM_cap_1_5_0[0|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|2]/vdd fgcell_amp_MiM_cap_1_5_0[0|2]/vsrc fgcell_amp_MiM_cap_1_5_0[0|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|2] fgcell_amp_MiM_cap_1_5_0[1|2]/vinj fgcell_amp_MiM_cap_1_5_0[1|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|2]/vdd fgcell_amp_MiM_cap_1_5_0[1|2]/vsrc fgcell_amp_MiM_cap_1_5_0[1|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|2] fgcell_amp_MiM_cap_1_5_0[2|2]/vinj fgcell_amp_MiM_cap_1_5_0[2|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|2]/vdd fgcell_amp_MiM_cap_1_5_0[2|2]/vsrc fgcell_amp_MiM_cap_1_5_0[2|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|2] fgcell_amp_MiM_cap_1_5_0[3|2]/vinj fgcell_amp_MiM_cap_1_5_0[3|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|2]/vdd fgcell_amp_MiM_cap_1_5_0[3|2]/vsrc fgcell_amp_MiM_cap_1_5_0[3|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|2] fgcell_amp_MiM_cap_1_5_0[4|2]/vinj fgcell_amp_MiM_cap_1_5_0[4|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|2]/vdd fgcell_amp_MiM_cap_1_5_0[4|2]/vsrc fgcell_amp_MiM_cap_1_5_0[4|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|2] fgcell_amp_MiM_cap_1_5_0[5|2]/vinj fgcell_amp_MiM_cap_1_5_0[5|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|2]/vdd fgcell_amp_MiM_cap_1_5_0[5|2]/vsrc fgcell_amp_MiM_cap_1_5_0[5|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|2] fgcell_amp_MiM_cap_1_5_0[6|2]/vinj fgcell_amp_MiM_cap_1_5_0[6|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|2]/vdd fgcell_amp_MiM_cap_1_5_0[6|2]/vsrc fgcell_amp_MiM_cap_1_5_0[6|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|2] fgcell_amp_MiM_cap_1_5_0[7|2]/vinj fgcell_amp_MiM_cap_1_5_0[7|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|2]/vdd fgcell_amp_MiM_cap_1_5_0[7|2]/vsrc fgcell_amp_MiM_cap_1_5_0[7|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|2] fgcell_amp_MiM_cap_1_5_0[8|2]/vinj fgcell_amp_MiM_cap_1_5_0[8|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|2]/vdd fgcell_amp_MiM_cap_1_5_0[8|2]/vsrc fgcell_amp_MiM_cap_1_5_0[8|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|2] fgcell_amp_MiM_cap_1_5_0[9|2]/vinj fgcell_amp_MiM_cap_1_5_0[9|2]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|2]/vdd fgcell_amp_MiM_cap_1_5_0[9|2]/vsrc fgcell_amp_MiM_cap_1_5_0[9|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|3] fgcell_amp_MiM_cap_1_5_0[0|3]/vinj fgcell_amp_MiM_cap_1_5_0[0|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|3]/vdd fgcell_amp_MiM_cap_1_5_0[0|3]/vsrc fgcell_amp_MiM_cap_1_5_0[0|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|3] fgcell_amp_MiM_cap_1_5_0[1|3]/vinj fgcell_amp_MiM_cap_1_5_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|3]/vdd fgcell_amp_MiM_cap_1_5_0[1|3]/vsrc fgcell_amp_MiM_cap_1_5_0[1|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|3] fgcell_amp_MiM_cap_1_5_0[2|3]/vinj fgcell_amp_MiM_cap_1_5_0[2|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|3]/vdd fgcell_amp_MiM_cap_1_5_0[2|3]/vsrc fgcell_amp_MiM_cap_1_5_0[2|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|3] fgcell_amp_MiM_cap_1_5_0[3|3]/vinj fgcell_amp_MiM_cap_1_5_0[3|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|3]/vdd fgcell_amp_MiM_cap_1_5_0[3|3]/vsrc fgcell_amp_MiM_cap_1_5_0[3|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|3] fgcell_amp_MiM_cap_1_5_0[4|3]/vinj fgcell_amp_MiM_cap_1_5_0[4|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|3]/vdd fgcell_amp_MiM_cap_1_5_0[4|3]/vsrc fgcell_amp_MiM_cap_1_5_0[4|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|3] fgcell_amp_MiM_cap_1_5_0[5|3]/vinj fgcell_amp_MiM_cap_1_5_0[5|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|3]/vdd fgcell_amp_MiM_cap_1_5_0[5|3]/vsrc fgcell_amp_MiM_cap_1_5_0[5|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|3] fgcell_amp_MiM_cap_1_5_0[6|3]/vinj fgcell_amp_MiM_cap_1_5_0[6|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|3]/vdd fgcell_amp_MiM_cap_1_5_0[6|3]/vsrc fgcell_amp_MiM_cap_1_5_0[6|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|3] fgcell_amp_MiM_cap_1_5_0[7|3]/vinj fgcell_amp_MiM_cap_1_5_0[7|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|3]/vdd fgcell_amp_MiM_cap_1_5_0[7|3]/vsrc fgcell_amp_MiM_cap_1_5_0[7|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|3] fgcell_amp_MiM_cap_1_5_0[8|3]/vinj fgcell_amp_MiM_cap_1_5_0[8|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|3]/vdd fgcell_amp_MiM_cap_1_5_0[8|3]/vsrc fgcell_amp_MiM_cap_1_5_0[8|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|3] fgcell_amp_MiM_cap_1_5_0[9|3]/vinj fgcell_amp_MiM_cap_1_5_0[9|3]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|3]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|3]/vdd fgcell_amp_MiM_cap_1_5_0[9|3]/vsrc fgcell_amp_MiM_cap_1_5_0[9|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|4] fgcell_amp_MiM_cap_1_5_0[0|4]/vinj fgcell_amp_MiM_cap_1_5_0[0|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|4]/vdd fgcell_amp_MiM_cap_1_5_0[0|4]/vsrc fgcell_amp_MiM_cap_1_5_0[0|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|4] fgcell_amp_MiM_cap_1_5_0[1|4]/vinj fgcell_amp_MiM_cap_1_5_0[1|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|4]/vdd fgcell_amp_MiM_cap_1_5_0[1|4]/vsrc fgcell_amp_MiM_cap_1_5_0[1|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|4] fgcell_amp_MiM_cap_1_5_0[2|4]/vinj fgcell_amp_MiM_cap_1_5_0[2|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|4]/vdd fgcell_amp_MiM_cap_1_5_0[2|4]/vsrc fgcell_amp_MiM_cap_1_5_0[2|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|4] fgcell_amp_MiM_cap_1_5_0[3|4]/vinj fgcell_amp_MiM_cap_1_5_0[3|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|4]/vdd fgcell_amp_MiM_cap_1_5_0[3|4]/vsrc fgcell_amp_MiM_cap_1_5_0[3|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|4] fgcell_amp_MiM_cap_1_5_0[4|4]/vinj fgcell_amp_MiM_cap_1_5_0[4|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|4]/vdd fgcell_amp_MiM_cap_1_5_0[4|4]/vsrc fgcell_amp_MiM_cap_1_5_0[4|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|4] fgcell_amp_MiM_cap_1_5_0[5|4]/vinj fgcell_amp_MiM_cap_1_5_0[5|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|4]/vdd fgcell_amp_MiM_cap_1_5_0[5|4]/vsrc fgcell_amp_MiM_cap_1_5_0[5|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|4] fgcell_amp_MiM_cap_1_5_0[6|4]/vinj fgcell_amp_MiM_cap_1_5_0[6|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|4]/vdd fgcell_amp_MiM_cap_1_5_0[6|4]/vsrc fgcell_amp_MiM_cap_1_5_0[6|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|4] fgcell_amp_MiM_cap_1_5_0[7|4]/vinj fgcell_amp_MiM_cap_1_5_0[7|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|4]/vdd fgcell_amp_MiM_cap_1_5_0[7|4]/vsrc fgcell_amp_MiM_cap_1_5_0[7|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|4] fgcell_amp_MiM_cap_1_5_0[8|4]/vinj fgcell_amp_MiM_cap_1_5_0[8|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|4]/vdd fgcell_amp_MiM_cap_1_5_0[8|4]/vsrc fgcell_amp_MiM_cap_1_5_0[8|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|4] fgcell_amp_MiM_cap_1_5_0[9|4]/vinj fgcell_amp_MiM_cap_1_5_0[9|4]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|4]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|4]/vdd fgcell_amp_MiM_cap_1_5_0[9|4]/vsrc fgcell_amp_MiM_cap_1_5_0[9|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|5] fgcell_amp_MiM_cap_1_5_0[0|5]/vinj fgcell_amp_MiM_cap_1_5_0[0|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|5]/vdd fgcell_amp_MiM_cap_1_5_0[0|5]/vsrc fgcell_amp_MiM_cap_1_5_0[0|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|5] fgcell_amp_MiM_cap_1_5_0[1|5]/vinj fgcell_amp_MiM_cap_1_5_0[1|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|5]/vdd fgcell_amp_MiM_cap_1_5_0[1|5]/vsrc fgcell_amp_MiM_cap_1_5_0[1|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|5] fgcell_amp_MiM_cap_1_5_0[2|5]/vinj fgcell_amp_MiM_cap_1_5_0[2|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|5]/vdd fgcell_amp_MiM_cap_1_5_0[2|5]/vsrc fgcell_amp_MiM_cap_1_5_0[2|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|5] fgcell_amp_MiM_cap_1_5_0[3|5]/vinj fgcell_amp_MiM_cap_1_5_0[3|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|5]/vdd fgcell_amp_MiM_cap_1_5_0[3|5]/vsrc fgcell_amp_MiM_cap_1_5_0[3|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|5] fgcell_amp_MiM_cap_1_5_0[4|5]/vinj fgcell_amp_MiM_cap_1_5_0[4|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|5]/vdd fgcell_amp_MiM_cap_1_5_0[4|5]/vsrc fgcell_amp_MiM_cap_1_5_0[4|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|5] fgcell_amp_MiM_cap_1_5_0[5|5]/vinj fgcell_amp_MiM_cap_1_5_0[5|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|5]/vdd fgcell_amp_MiM_cap_1_5_0[5|5]/vsrc fgcell_amp_MiM_cap_1_5_0[5|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|5] fgcell_amp_MiM_cap_1_5_0[6|5]/vinj fgcell_amp_MiM_cap_1_5_0[6|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|5]/vdd fgcell_amp_MiM_cap_1_5_0[6|5]/vsrc fgcell_amp_MiM_cap_1_5_0[6|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|5] fgcell_amp_MiM_cap_1_5_0[7|5]/vinj fgcell_amp_MiM_cap_1_5_0[7|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|5]/vdd fgcell_amp_MiM_cap_1_5_0[7|5]/vsrc fgcell_amp_MiM_cap_1_5_0[7|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|5] fgcell_amp_MiM_cap_1_5_0[8|5]/vinj fgcell_amp_MiM_cap_1_5_0[8|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|5]/vdd fgcell_amp_MiM_cap_1_5_0[8|5]/vsrc fgcell_amp_MiM_cap_1_5_0[8|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|5] fgcell_amp_MiM_cap_1_5_0[9|5]/vinj fgcell_amp_MiM_cap_1_5_0[9|5]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|5]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|5]/vdd fgcell_amp_MiM_cap_1_5_0[9|5]/vsrc fgcell_amp_MiM_cap_1_5_0[9|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|6] fgcell_amp_MiM_cap_1_5_0[0|6]/vinj fgcell_amp_MiM_cap_1_5_0[0|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|6]/vdd fgcell_amp_MiM_cap_1_5_0[0|6]/vsrc fgcell_amp_MiM_cap_1_5_0[0|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|6] fgcell_amp_MiM_cap_1_5_0[1|6]/vinj fgcell_amp_MiM_cap_1_5_0[1|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|6]/vdd fgcell_amp_MiM_cap_1_5_0[1|6]/vsrc fgcell_amp_MiM_cap_1_5_0[1|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|6] fgcell_amp_MiM_cap_1_5_0[2|6]/vinj fgcell_amp_MiM_cap_1_5_0[2|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|6]/vdd fgcell_amp_MiM_cap_1_5_0[2|6]/vsrc fgcell_amp_MiM_cap_1_5_0[2|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|6] fgcell_amp_MiM_cap_1_5_0[3|6]/vinj fgcell_amp_MiM_cap_1_5_0[3|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|6]/vdd fgcell_amp_MiM_cap_1_5_0[3|6]/vsrc fgcell_amp_MiM_cap_1_5_0[3|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|6] fgcell_amp_MiM_cap_1_5_0[4|6]/vinj fgcell_amp_MiM_cap_1_5_0[4|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|6]/vdd fgcell_amp_MiM_cap_1_5_0[4|6]/vsrc fgcell_amp_MiM_cap_1_5_0[4|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|6] fgcell_amp_MiM_cap_1_5_0[5|6]/vinj fgcell_amp_MiM_cap_1_5_0[5|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|6]/vdd fgcell_amp_MiM_cap_1_5_0[5|6]/vsrc fgcell_amp_MiM_cap_1_5_0[5|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|6] fgcell_amp_MiM_cap_1_5_0[6|6]/vinj fgcell_amp_MiM_cap_1_5_0[6|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|6]/vdd fgcell_amp_MiM_cap_1_5_0[6|6]/vsrc fgcell_amp_MiM_cap_1_5_0[6|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|6] fgcell_amp_MiM_cap_1_5_0[7|6]/vinj fgcell_amp_MiM_cap_1_5_0[7|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|6]/vdd fgcell_amp_MiM_cap_1_5_0[7|6]/vsrc fgcell_amp_MiM_cap_1_5_0[7|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|6] fgcell_amp_MiM_cap_1_5_0[8|6]/vinj fgcell_amp_MiM_cap_1_5_0[8|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|6]/vdd fgcell_amp_MiM_cap_1_5_0[8|6]/vsrc fgcell_amp_MiM_cap_1_5_0[8|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|6] fgcell_amp_MiM_cap_1_5_0[9|6]/vinj fgcell_amp_MiM_cap_1_5_0[9|6]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|6]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|6]/vdd fgcell_amp_MiM_cap_1_5_0[9|6]/vsrc fgcell_amp_MiM_cap_1_5_0[9|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|7] fgcell_amp_MiM_cap_1_5_0[0|7]/vinj fgcell_amp_MiM_cap_1_5_0[0|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|7]/vdd fgcell_amp_MiM_cap_1_5_0[0|7]/vsrc fgcell_amp_MiM_cap_1_5_0[0|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|7] fgcell_amp_MiM_cap_1_5_0[1|7]/vinj fgcell_amp_MiM_cap_1_5_0[1|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|7]/vdd fgcell_amp_MiM_cap_1_5_0[1|7]/vsrc fgcell_amp_MiM_cap_1_5_0[1|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|7] fgcell_amp_MiM_cap_1_5_0[2|7]/vinj fgcell_amp_MiM_cap_1_5_0[2|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|7]/vdd fgcell_amp_MiM_cap_1_5_0[2|7]/vsrc fgcell_amp_MiM_cap_1_5_0[2|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|7] fgcell_amp_MiM_cap_1_5_0[3|7]/vinj fgcell_amp_MiM_cap_1_5_0[3|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|7]/vdd fgcell_amp_MiM_cap_1_5_0[3|7]/vsrc fgcell_amp_MiM_cap_1_5_0[3|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|7] fgcell_amp_MiM_cap_1_5_0[4|7]/vinj fgcell_amp_MiM_cap_1_5_0[4|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|7]/vdd fgcell_amp_MiM_cap_1_5_0[4|7]/vsrc fgcell_amp_MiM_cap_1_5_0[4|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|7] fgcell_amp_MiM_cap_1_5_0[5|7]/vinj fgcell_amp_MiM_cap_1_5_0[5|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|7]/vdd fgcell_amp_MiM_cap_1_5_0[5|7]/vsrc fgcell_amp_MiM_cap_1_5_0[5|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|7] fgcell_amp_MiM_cap_1_5_0[6|7]/vinj fgcell_amp_MiM_cap_1_5_0[6|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|7]/vdd fgcell_amp_MiM_cap_1_5_0[6|7]/vsrc fgcell_amp_MiM_cap_1_5_0[6|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|7] fgcell_amp_MiM_cap_1_5_0[7|7]/vinj fgcell_amp_MiM_cap_1_5_0[7|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|7]/vdd fgcell_amp_MiM_cap_1_5_0[7|7]/vsrc fgcell_amp_MiM_cap_1_5_0[7|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|7] fgcell_amp_MiM_cap_1_5_0[8|7]/vinj fgcell_amp_MiM_cap_1_5_0[8|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|7]/vdd fgcell_amp_MiM_cap_1_5_0[8|7]/vsrc fgcell_amp_MiM_cap_1_5_0[8|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|7] fgcell_amp_MiM_cap_1_5_0[9|7]/vinj fgcell_amp_MiM_cap_1_5_0[9|7]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|7]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|7]/vdd fgcell_amp_MiM_cap_1_5_0[9|7]/vsrc fgcell_amp_MiM_cap_1_5_0[9|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|8] fgcell_amp_MiM_cap_1_5_0[0|8]/vinj fgcell_amp_MiM_cap_1_5_0[0|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|8]/vdd fgcell_amp_MiM_cap_1_5_0[0|8]/vsrc fgcell_amp_MiM_cap_1_5_0[0|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|8] fgcell_amp_MiM_cap_1_5_0[1|8]/vinj fgcell_amp_MiM_cap_1_5_0[1|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|8]/vdd fgcell_amp_MiM_cap_1_5_0[1|8]/vsrc fgcell_amp_MiM_cap_1_5_0[1|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|8] fgcell_amp_MiM_cap_1_5_0[2|8]/vinj fgcell_amp_MiM_cap_1_5_0[2|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|8]/vdd fgcell_amp_MiM_cap_1_5_0[2|8]/vsrc fgcell_amp_MiM_cap_1_5_0[2|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|8] fgcell_amp_MiM_cap_1_5_0[3|8]/vinj fgcell_amp_MiM_cap_1_5_0[3|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|8]/vdd fgcell_amp_MiM_cap_1_5_0[3|8]/vsrc fgcell_amp_MiM_cap_1_5_0[3|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|8] fgcell_amp_MiM_cap_1_5_0[4|8]/vinj fgcell_amp_MiM_cap_1_5_0[4|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|8]/vdd fgcell_amp_MiM_cap_1_5_0[4|8]/vsrc fgcell_amp_MiM_cap_1_5_0[4|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|8] fgcell_amp_MiM_cap_1_5_0[5|8]/vinj fgcell_amp_MiM_cap_1_5_0[5|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|8]/vdd fgcell_amp_MiM_cap_1_5_0[5|8]/vsrc fgcell_amp_MiM_cap_1_5_0[5|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|8] fgcell_amp_MiM_cap_1_5_0[6|8]/vinj fgcell_amp_MiM_cap_1_5_0[6|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|8]/vdd fgcell_amp_MiM_cap_1_5_0[6|8]/vsrc fgcell_amp_MiM_cap_1_5_0[6|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|8] fgcell_amp_MiM_cap_1_5_0[7|8]/vinj fgcell_amp_MiM_cap_1_5_0[7|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|8]/vdd fgcell_amp_MiM_cap_1_5_0[7|8]/vsrc fgcell_amp_MiM_cap_1_5_0[7|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|8] fgcell_amp_MiM_cap_1_5_0[8|8]/vinj fgcell_amp_MiM_cap_1_5_0[8|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|8]/vdd fgcell_amp_MiM_cap_1_5_0[8|8]/vsrc fgcell_amp_MiM_cap_1_5_0[8|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|8] fgcell_amp_MiM_cap_1_5_0[9|8]/vinj fgcell_amp_MiM_cap_1_5_0[9|8]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|8]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|8]/vdd fgcell_amp_MiM_cap_1_5_0[9|8]/vsrc fgcell_amp_MiM_cap_1_5_0[9|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[0|9] fgcell_amp_MiM_cap_1_5_0[0|9]/vinj fgcell_amp_MiM_cap_1_5_0[0|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[0|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[0|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[0|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[0|9]/vdd fgcell_amp_MiM_cap_1_5_0[0|9]/vsrc fgcell_amp_MiM_cap_1_5_0[0|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[1|9] fgcell_amp_MiM_cap_1_5_0[1|9]/vinj fgcell_amp_MiM_cap_1_5_0[1|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[1|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[1|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[1|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[1|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[1|9]/vdd fgcell_amp_MiM_cap_1_5_0[1|9]/vsrc fgcell_amp_MiM_cap_1_5_0[1|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[2|9] fgcell_amp_MiM_cap_1_5_0[2|9]/vinj fgcell_amp_MiM_cap_1_5_0[2|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[2|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[2|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[2|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[2|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[2|9]/vdd fgcell_amp_MiM_cap_1_5_0[2|9]/vsrc fgcell_amp_MiM_cap_1_5_0[2|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[3|9] fgcell_amp_MiM_cap_1_5_0[3|9]/vinj fgcell_amp_MiM_cap_1_5_0[3|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[3|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[3|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[3|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[3|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[3|9]/vdd fgcell_amp_MiM_cap_1_5_0[3|9]/vsrc fgcell_amp_MiM_cap_1_5_0[3|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[4|9] fgcell_amp_MiM_cap_1_5_0[4|9]/vinj fgcell_amp_MiM_cap_1_5_0[4|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[4|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[4|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[4|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[4|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[4|9]/vdd fgcell_amp_MiM_cap_1_5_0[4|9]/vsrc fgcell_amp_MiM_cap_1_5_0[4|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[5|9] fgcell_amp_MiM_cap_1_5_0[5|9]/vinj fgcell_amp_MiM_cap_1_5_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[5|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[5|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[5|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[5|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[5|9]/vdd fgcell_amp_MiM_cap_1_5_0[5|9]/vsrc fgcell_amp_MiM_cap_1_5_0[5|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[6|9] fgcell_amp_MiM_cap_1_5_0[6|9]/vinj fgcell_amp_MiM_cap_1_5_0[6|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[6|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[6|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[6|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[6|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[6|9]/vdd fgcell_amp_MiM_cap_1_5_0[6|9]/vsrc fgcell_amp_MiM_cap_1_5_0[6|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[7|9] fgcell_amp_MiM_cap_1_5_0[7|9]/vinj fgcell_amp_MiM_cap_1_5_0[7|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[7|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[7|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[7|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[7|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[7|9]/vdd fgcell_amp_MiM_cap_1_5_0[7|9]/vsrc fgcell_amp_MiM_cap_1_5_0[7|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[8|9] fgcell_amp_MiM_cap_1_5_0[8|9]/vinj fgcell_amp_MiM_cap_1_5_0[8|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[8|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[8|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[8|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[8|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[8|9]/vdd fgcell_amp_MiM_cap_1_5_0[8|9]/vsrc fgcell_amp_MiM_cap_1_5_0[8|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
Xfgcell_amp_MiM_cap_1_5_0[9|9] fgcell_amp_MiM_cap_1_5_0[9|9]/vinj fgcell_amp_MiM_cap_1_5_0[9|9]/vtun
+ fgcell_amp_MiM_cap_1_5_0[9|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_5_0[9|9]/row_en
+ fgcell_amp_MiM_cap_1_5_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_5_0[9|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_5_0[9|9]/vdd fgcell_amp_MiM_cap_1_5_0[9|9]/vsrc fgcell_amp_MiM_cap_1_5_0[9|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_5
.ends

.subckt lsi1v8o5v0 in out_b out vdd_l vdd_h vss
X0 vdd_l in in_b vdd_l sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X1 vss t1 out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X2 out_b out vdd_h vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X3 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=1.305 ps=14.22 w=0.5 l=0.5
X4 vdd_h out out_b vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X5 out_b out vdd_h vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X6 vss in in_b vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X7 vdd_h out out_b vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X8 in_bb in_b vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X9 vdd_h t1 out vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X10 out t1 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X11 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=0.5
X12 vdd_h t1 out vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X13 in_bb in_b vdd_l vdd_l sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X14 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=0.5
X15 vdd_h t1 t2 vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X16 out t1 vdd_h vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X17 t1 in_bb vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X18 out t1 vdd_h vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X19 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=0.5
X20 t1 t2 vdd_h vdd_h sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X21 out_b out vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
X22 vss in_b t2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X23 vss out out_b vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.5
.ends

.subckt fgcell_amp_MiM_cap_1_10 vinj vtun x1/tg5v0_0/vout row_en x1/x1/vctrl x1/x2/vb
+ vdd vsrc row_en_b VGND
Xx1 vtun x1/tg5v0_0/vout vdd x1/x2/v1 row_en vsrc x1/x1/vctrl row_en_b VGND vinj x1/x2/vb
+ fgcell_amp
X0 x1/x2/v1 VGND sky130_fd_pr__cap_mim_m3_1 l=1 w=10
.ends

.subckt array_core_block2 fgcell_amp_MiM_cap_1_10_0[9|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[3|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|2]/vsrc fgcell_amp_MiM_cap_1_10_0[6|5]/row_en_b fgcell_amp_MiM_cap_1_10_0[6|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|7]/vsrc fgcell_amp_MiM_cap_1_10_0[9|9]/vsrc fgcell_amp_MiM_cap_1_10_0[4|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|8]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[7|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[9|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[6|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[1|5]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[6|0]/vtun fgcell_amp_MiM_cap_1_10_0[2|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|5]/vtun fgcell_amp_MiM_cap_1_10_0[4|3]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[1|8]/vsrc fgcell_amp_MiM_cap_1_10_0[8|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[7|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[8|5]/vdd fgcell_amp_MiM_cap_1_10_0[6|4]/vinj
+ fgcell_amp_MiM_cap_1_10_0[6|1]/vtun fgcell_amp_MiM_cap_1_10_0[6|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|6]/vtun fgcell_amp_MiM_cap_1_10_0[4|4]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[3|8]/vinj fgcell_amp_MiM_cap_1_10_0[1|9]/vsrc fgcell_amp_MiM_cap_1_10_0[9|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|5]/vinj fgcell_amp_MiM_cap_1_10_0[9|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[7|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[3|7]/vtun fgcell_amp_MiM_cap_1_10_0[7|0]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[4|5]/vsrc fgcell_amp_MiM_cap_1_10_0[7|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[8|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[2|3]/vdd fgcell_amp_MiM_cap_1_10_0[1|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[8|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|9]/vinj fgcell_amp_MiM_cap_1_10_0[2|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[6|6]/vinj
+ fgcell_amp_MiM_cap_1_10_0[6|3]/vtun fgcell_amp_MiM_cap_1_10_0[1|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|1]/vsrc fgcell_amp_MiM_cap_1_10_0[3|8]/vtun fgcell_amp_MiM_cap_1_10_0[0|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[8|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[6|7]/vinj fgcell_amp_MiM_cap_1_10_0[6|4]/vtun fgcell_amp_MiM_cap_1_10_0[9|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|2]/vsrc fgcell_amp_MiM_cap_1_10_0[4|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[4|7]/vsrc fgcell_amp_MiM_cap_1_10_0[0|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[4|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|0]/vtun fgcell_amp_MiM_cap_1_10_0[6|8]/vinj fgcell_amp_MiM_cap_1_10_0[8|6]/vdd
+ fgcell_amp_MiM_cap_1_10_0[6|5]/vtun fgcell_amp_MiM_cap_1_10_0[7|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[7|3]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[7|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|1]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[4|8]/vsrc fgcell_amp_MiM_cap_1_10_0[0|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|4]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|7]/vdd fgcell_amp_MiM_cap_1_10_0[7|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|6]/vdd fgcell_amp_MiM_cap_1_10_0[9|1]/vtun fgcell_amp_MiM_cap_1_10_0[3|1]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[0|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[6|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[0|2]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|9]/vtun fgcell_amp_MiM_cap_1_10_0[0|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|4]/row_en_b fgcell_amp_MiM_cap_1_10_0[7|4]/vsrc fgcell_amp_MiM_cap_1_10_0[4|9]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[3|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[9|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|4]/vdd fgcell_amp_MiM_cap_1_10_0[1|2]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|5]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[6|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|2]/vdd
+ fgcell_amp_MiM_cap_1_10_0[3|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[9|3]/vtun fgcell_amp_MiM_cap_1_10_0[2|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|8]/vtun fgcell_amp_MiM_cap_1_10_0[9|9]/vdd fgcell_amp_MiM_cap_1_10_0[8|5]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[6|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|8]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[6|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|0]/vinj fgcell_amp_MiM_cap_1_10_0[3|5]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|8]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|4]/vtun fgcell_amp_MiM_cap_1_10_0[3|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|0]/vsrc fgcell_amp_MiM_cap_1_10_0[1|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[7|7]/vsrc fgcell_amp_MiM_cap_1_10_0[7|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[4|1]/vinj fgcell_amp_MiM_cap_1_10_0[9|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[9|5]/vtun fgcell_amp_MiM_cap_1_10_0[4|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|1]/vsrc fgcell_amp_MiM_cap_1_10_0[2|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[7|8]/vsrc fgcell_amp_MiM_cap_1_10_0[6|2]/vdd fgcell_amp_MiM_cap_1_10_0[1|0]/vinj
+ fgcell_amp_MiM_cap_1_10_0[5|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|7]/vdd
+ fgcell_amp_MiM_cap_1_10_0[4|2]/vinj fgcell_amp_MiM_cap_1_10_0[6|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|5]/vdd
+ fgcell_amp_MiM_cap_1_10_0[8|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|2]/vsrc fgcell_amp_MiM_cap_1_10_0[5|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[7|9]/vsrc fgcell_amp_MiM_cap_1_10_0[6|6]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[3|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[7|0]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|3]/vinj fgcell_amp_MiM_cap_1_10_0[4|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|3]/vdd fgcell_amp_MiM_cap_1_10_0[7|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[1|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|7]/vtun fgcell_amp_MiM_cap_1_10_0[5|1]/vdd
+ fgcell_amp_MiM_cap_1_10_0[6|2]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|3]/vsrc fgcell_amp_MiM_cap_1_10_0[1|1]/vinj
+ fgcell_amp_MiM_cap_1_10_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|0]/vinj fgcell_amp_MiM_cap_1_10_0[4|4]/vinj fgcell_amp_MiM_cap_1_10_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|1]/vdd fgcell_amp_MiM_cap_1_10_0[8|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[4|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|8]/vtun fgcell_amp_MiM_cap_1_10_0[2|4]/vsrc fgcell_amp_MiM_cap_1_10_0[2|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|2]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[4|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|0]/vtun fgcell_amp_MiM_cap_1_10_0[1|2]/vinj fgcell_amp_MiM_cap_1_10_0[3|7]/vdd
+ fgcell_amp_MiM_cap_1_10_0[4|5]/vinj fgcell_amp_MiM_cap_1_10_0[9|6]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[4|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|0]/vsrc fgcell_amp_MiM_cap_1_10_0[7|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[8|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|5]/vsrc fgcell_amp_MiM_cap_1_10_0[7|6]/vdd fgcell_amp_MiM_cap_1_10_0[9|1]/vinj
+ fgcell_amp_MiM_cap_1_10_0[0|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[4|6]/vinj fgcell_amp_MiM_cap_1_10_0[5|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[5|1]/vsrc fgcell_amp_MiM_cap_1_10_0[2|6]/vdd fgcell_amp_MiM_cap_1_10_0[0|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[9|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|1]/vtun fgcell_amp_MiM_cap_1_10_0[1|3]/vinj fgcell_amp_MiM_cap_1_10_0[0|1]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[4|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|7]/vinj fgcell_amp_MiM_cap_1_10_0[4|4]/vtun fgcell_amp_MiM_cap_1_10_0[9|2]/vinj
+ fgcell_amp_MiM_cap_1_10_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[5|2]/vsrc fgcell_amp_MiM_cap_1_10_0[1|4]/vdd fgcell_amp_MiM_cap_1_10_0[2|7]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[7|3]/vdd fgcell_amp_MiM_cap_1_10_0[9|0]/vdd fgcell_amp_MiM_cap_1_10_0[3|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|9]/vtun fgcell_amp_MiM_cap_1_10_0[1|7]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[7|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|8]/vinj fgcell_amp_MiM_cap_1_10_0[1|2]/vtun fgcell_amp_MiM_cap_1_10_0[4|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|2]/vdd fgcell_amp_MiM_cap_1_10_0[1|4]/vinj fgcell_amp_MiM_cap_1_10_0[6|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[4|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|3]/vsrc fgcell_amp_MiM_cap_1_10_0[2|8]/vsrc fgcell_amp_MiM_cap_1_10_0[7|8]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[8|9]/vdd fgcell_amp_MiM_cap_1_10_0[8|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|3]/vinj
+ fgcell_amp_MiM_cap_1_10_0[6|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|5]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[7|1]/vtun fgcell_amp_MiM_cap_1_10_0[2|8]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|9]/vinj fgcell_amp_MiM_cap_1_10_0[4|6]/vtun fgcell_amp_MiM_cap_1_10_0[3|2]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|4]/vsrc fgcell_amp_MiM_cap_1_10_0[9|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|5]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|9]/vsrc fgcell_amp_MiM_cap_1_10_0[5|2]/vdd
+ fgcell_amp_MiM_cap_1_10_0[2|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|5]/vinj fgcell_amp_MiM_cap_1_10_0[8|7]/vdd fgcell_amp_MiM_cap_1_10_0[9|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|7]/vtun fgcell_amp_MiM_cap_1_10_0[8|0]/vsrc fgcell_amp_MiM_cap_1_10_0[2|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|2]/vtun fgcell_amp_MiM_cap_1_10_0[2|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|5]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[9|4]/vinj fgcell_amp_MiM_cap_1_10_0[8|3]/row_en fgcell_amp_MiM_cap_1_10_0[6|5]/vdd
+ fgcell_amp_MiM_cap_1_10_0[5|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|8]/vdd fgcell_amp_MiM_cap_1_10_0[7|6]/vinj fgcell_amp_MiM_cap_1_10_0[4|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|3]/vtun fgcell_amp_MiM_cap_1_10_0[4|9]/row_en fgcell_amp_MiM_cap_1_10_0[8|1]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[4|8]/vtun fgcell_amp_MiM_cap_1_10_0[5|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[3|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|6]/vsrc fgcell_amp_MiM_cap_1_10_0[1|5]/vdd
+ fgcell_amp_MiM_cap_1_10_0[1|4]/vtun fgcell_amp_MiM_cap_1_10_0[8|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|6]/vinj
+ fgcell_amp_MiM_cap_1_10_0[2|6]/vsrc fgcell_amp_MiM_cap_1_10_0[5|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[8|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|1]/vdd fgcell_amp_MiM_cap_1_10_0[6|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|9]/vdd
+ fgcell_amp_MiM_cap_1_10_0[9|5]/vinj fgcell_amp_MiM_cap_1_10_0[1|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[8|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|4]/vtun fgcell_amp_MiM_cap_1_10_0[7|7]/vinj
+ fgcell_amp_MiM_cap_1_10_0[3|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[5|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|0]/vsrc fgcell_amp_MiM_cap_1_10_0[4|9]/vtun fgcell_amp_MiM_cap_1_10_0[8|2]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[0|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[8|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[4|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|7]/vsrc fgcell_amp_MiM_cap_1_10_0[1|3]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[4|1]/vdd fgcell_amp_MiM_cap_1_10_0[1|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[7|5]/row_en fgcell_amp_MiM_cap_1_10_0[8|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[2|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[1|5]/vtun fgcell_amp_MiM_cap_1_10_0[7|8]/vinj fgcell_amp_MiM_cap_1_10_0[6|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|5]/vtun fgcell_amp_MiM_cap_1_10_0[1|7]/vinj fgcell_amp_MiM_cap_1_10_0[2|7]/vdd
+ fgcell_amp_MiM_cap_1_10_0[0|5]/row_en fgcell_amp_MiM_cap_1_10_0[0|1]/vsrc fgcell_amp_MiM_cap_1_10_0[8|3]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[5|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|8]/vsrc fgcell_amp_MiM_cap_1_10_0[2|0]/vinj
+ fgcell_amp_MiM_cap_1_10_0[7|0]/row_en fgcell_amp_MiM_cap_1_10_0[9|6]/vinj fgcell_amp_MiM_cap_1_10_0[4|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|0]/row_en fgcell_amp_MiM_cap_1_10_0[1|0]/vdd fgcell_amp_MiM_cap_1_10_0[7|9]/vinj
+ fgcell_amp_MiM_cap_1_10_0[7|6]/vtun fgcell_amp_MiM_cap_1_10_0[3|6]/row_en fgcell_amp_MiM_cap_1_10_0[7|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|2]/vsrc fgcell_amp_MiM_cap_1_10_0[8|4]/vsrc fgcell_amp_MiM_cap_1_10_0[4|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|9]/vsrc fgcell_amp_MiM_cap_1_10_0[6|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[9|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|6]/vtun fgcell_amp_MiM_cap_1_10_0[6|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|8]/vinj
+ fgcell_amp_MiM_cap_1_10_0[6|6]/vdd fgcell_amp_MiM_cap_1_10_0[3|1]/row_en fgcell_amp_MiM_cap_1_10_0[7|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[6|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|0]/vtun fgcell_amp_MiM_cap_1_10_0[2|1]/vinj
+ fgcell_amp_MiM_cap_1_10_0[0|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|7]/vtun fgcell_amp_MiM_cap_1_10_0[6|7]/row_en fgcell_amp_MiM_cap_1_10_0[0|3]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[8|5]/vsrc fgcell_amp_MiM_cap_1_10_0[9|7]/vinj fgcell_amp_MiM_cap_1_10_0[1|7]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|6]/vdd fgcell_amp_MiM_cap_1_10_0[6|3]/vdd
+ fgcell_amp_MiM_cap_1_10_0[0|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[9|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|4]/vdd fgcell_amp_MiM_cap_1_10_0[6|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|2]/vdd fgcell_amp_MiM_cap_1_10_0[9|8]/vdd fgcell_amp_MiM_cap_1_10_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|8]/vtun fgcell_amp_MiM_cap_1_10_0[9|7]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[1|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|4]/vsrc fgcell_amp_MiM_cap_1_10_0[9|8]/row_en fgcell_amp_MiM_cap_1_10_0[8|6]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[1|9]/vinj fgcell_amp_MiM_cap_1_10_0[0|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|8]/row_en fgcell_amp_MiM_cap_1_10_0[5|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|2]/vinj fgcell_amp_MiM_cap_1_10_0[3|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|6]/vtun fgcell_amp_MiM_cap_1_10_0[5|0]/vinj fgcell_amp_MiM_cap_1_10_0[9|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|9]/vdd fgcell_amp_MiM_cap_1_10_0[8|0]/vdd fgcell_amp_MiM_cap_1_10_0[9|8]/vinj
+ fgcell_amp_MiM_cap_1_10_0[8|9]/row_en fgcell_amp_MiM_cap_1_10_0[3|0]/vsrc fgcell_amp_MiM_cap_1_10_0[6|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|3]/row_en fgcell_amp_MiM_cap_1_10_0[7|9]/vtun fgcell_amp_MiM_cap_1_10_0[0|5]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[8|7]/vsrc fgcell_amp_MiM_cap_1_10_0[9|8]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|3]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|9]/row_en fgcell_amp_MiM_cap_1_10_0[3|0]/vdd
+ fgcell_amp_MiM_cap_1_10_0[8|4]/row_en fgcell_amp_MiM_cap_1_10_0[7|5]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|1]/vinj
+ fgcell_amp_MiM_cap_1_10_0[4|2]/vdd fgcell_amp_MiM_cap_1_10_0[6|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|8]/vtun fgcell_amp_MiM_cap_1_10_0[7|9]/vdd fgcell_amp_MiM_cap_1_10_0[2|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|4]/row_en fgcell_amp_MiM_cap_1_10_0[4|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|1]/vsrc fgcell_amp_MiM_cap_1_10_0[7|7]/vdd fgcell_amp_MiM_cap_1_10_0[9|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|2]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|4]/row_en fgcell_amp_MiM_cap_1_10_0[2|3]/vinj
+ fgcell_amp_MiM_cap_1_10_0[2|5]/row_en_b fgcell_amp_MiM_cap_1_10_0[8|8]/vsrc fgcell_amp_MiM_cap_1_10_0[9|9]/vinj
+ fgcell_amp_MiM_cap_1_10_0[2|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[4|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[2|9]/vdd fgcell_amp_MiM_cap_1_10_0[0|3]/vdd fgcell_amp_MiM_cap_1_10_0[0|2]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|2]/vinj
+ fgcell_amp_MiM_cap_1_10_0[2|4]/vtun fgcell_amp_MiM_cap_1_10_0[4|5]/row_en fgcell_amp_MiM_cap_1_10_0[1|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|8]/vdd fgcell_amp_MiM_cap_1_10_0[2|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[3|2]/vsrc fgcell_amp_MiM_cap_1_10_0[8|5]/row_en fgcell_amp_MiM_cap_1_10_0[4|3]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|7]/vsrc fgcell_amp_MiM_cap_1_10_0[8|9]/vsrc fgcell_amp_MiM_cap_1_10_0[6|3]/vinj
+ fgcell_amp_MiM_cap_1_10_0[1|9]/vtun fgcell_amp_MiM_cap_1_10_0[1|5]/row_en fgcell_amp_MiM_cap_1_10_0[4|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|2]/vtun fgcell_amp_MiM_cap_1_10_0[5|3]/vinj fgcell_amp_MiM_cap_1_10_0[8|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|0]/vtun fgcell_amp_MiM_cap_1_10_0[2|4]/vinj fgcell_amp_MiM_cap_1_10_0[5|5]/vdd
+ fgcell_amp_MiM_cap_1_10_0[2|5]/vtun fgcell_amp_MiM_cap_1_10_0[9|3]/vdd fgcell_amp_MiM_cap_1_10_0[7|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|3]/vsrc fgcell_amp_MiM_cap_1_10_0[1|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|8]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[1|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[0|6]/row_en fgcell_amp_MiM_cap_1_10_0[7|9]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[4|6]/row_en fgcell_amp_MiM_cap_1_10_0[0|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[0|5]/vdd
+ fgcell_amp_MiM_cap_1_10_0[7|1]/row_en fgcell_amp_MiM_cap_1_10_0[8|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[5|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[6|2]/vtun fgcell_amp_MiM_cap_1_10_0[5|4]/vinj fgcell_amp_MiM_cap_1_10_0[5|6]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[5|1]/vtun fgcell_amp_MiM_cap_1_10_0[8|1]/vdd fgcell_amp_MiM_cap_1_10_0[0|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|9]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[3|4]/vsrc fgcell_amp_MiM_cap_1_10_0[4|1]/row_en fgcell_amp_MiM_cap_1_10_0[0|9]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[1|7]/vdd fgcell_amp_MiM_cap_1_10_0[3|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[5|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[2|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|7]/row_en fgcell_amp_MiM_cap_1_10_0[2|5]/vinj
+ fgcell_amp_MiM_cap_1_10_0[7|4]/vdd fgcell_amp_MiM_cap_1_10_0[0|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[1|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[9|9]/vtun fgcell_amp_MiM_cap_1_10_0[8|0]/vinj
+ fgcell_amp_MiM_cap_1_10_0[7|7]/row_en fgcell_amp_MiM_cap_1_10_0[1|0]/row_en_b fgcell_amp_MiM_cap_1_10_0[8|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[3|1]/vdd fgcell_amp_MiM_cap_1_10_0[5|5]/vinj fgcell_amp_MiM_cap_1_10_0[5|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|7]/row_en fgcell_amp_MiM_cap_1_10_0[6|0]/vsrc fgcell_amp_MiM_cap_1_10_0[3|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|7]/vtun fgcell_amp_MiM_cap_1_10_0[0|0]/vdd fgcell_amp_MiM_cap_1_10_0[1|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|5]/vsrc fgcell_amp_MiM_cap_1_10_0[7|2]/row_en fgcell_amp_MiM_cap_1_10_0[3|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|5]/vdd fgcell_amp_MiM_cap_1_10_0[6|8]/row_en fgcell_amp_MiM_cap_1_10_0[4|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|2]/row_en fgcell_amp_MiM_cap_1_10_0[2|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[8|1]/vinj
+ fgcell_amp_MiM_cap_1_10_0[5|6]/vinj fgcell_amp_MiM_cap_1_10_0[5|3]/vtun fgcell_amp_MiM_cap_1_10_0[6|8]/vdd
+ fgcell_amp_MiM_cap_1_10_0[3|8]/row_en fgcell_amp_MiM_cap_1_10_0[2|8]/vtun fgcell_amp_MiM_cap_1_10_0[6|1]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[6|3]/row_en fgcell_amp_MiM_cap_1_10_0[5|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|6]/vinj
+ fgcell_amp_MiM_cap_1_10_0[4|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|6]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[4|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[7|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[8|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|9]/row_en fgcell_amp_MiM_cap_1_10_0[5|3]/vdd
+ fgcell_amp_MiM_cap_1_10_0[3|3]/row_en fgcell_amp_MiM_cap_1_10_0[3|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[8|2]/vinj
+ fgcell_amp_MiM_cap_1_10_0[9|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|9]/row_en fgcell_amp_MiM_cap_1_10_0[5|7]/vinj
+ fgcell_amp_MiM_cap_1_10_0[0|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[5|4]/vtun fgcell_amp_MiM_cap_1_10_0[5|6]/vdd fgcell_amp_MiM_cap_1_10_0[8|8]/vdd
+ fgcell_amp_MiM_cap_1_10_0[6|2]/vsrc fgcell_amp_MiM_cap_1_10_0[6|9]/row_en fgcell_amp_MiM_cap_1_10_0[6|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[9|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|4]/vdd fgcell_amp_MiM_cap_1_10_0[3|7]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|4]/row_en fgcell_amp_MiM_cap_1_10_0[7|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[3|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|7]/vsrc fgcell_amp_MiM_cap_1_10_0[7|6]/vsrc fgcell_amp_MiM_cap_1_10_0[4|1]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[2|4]/row_en fgcell_amp_MiM_cap_1_10_0[5|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[1|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[0|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|1]/vinj fgcell_amp_MiM_cap_1_10_0[4|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[0|6]/vdd
+ fgcell_amp_MiM_cap_1_10_0[2|7]/vinj fgcell_amp_MiM_cap_1_10_0[8|3]/vinj fgcell_amp_MiM_cap_1_10_0[8|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[4|4]/vdd fgcell_amp_MiM_cap_1_10_0[5|8]/vinj fgcell_amp_MiM_cap_1_10_0[3|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[5|5]/vtun fgcell_amp_MiM_cap_1_10_0[4|9]/vdd fgcell_amp_MiM_cap_1_10_0[6|3]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[8|2]/vdd fgcell_amp_MiM_cap_1_10_0[7|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|8]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[6|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|5]/row_en fgcell_amp_MiM_cap_1_10_0[3|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|5]/row_en fgcell_amp_MiM_cap_1_10_0[5|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[0|2]/vinj
+ fgcell_amp_MiM_cap_1_10_0[8|4]/vinj fgcell_amp_MiM_cap_1_10_0[0|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|2]/vdd fgcell_amp_MiM_cap_1_10_0[5|9]/vinj fgcell_amp_MiM_cap_1_10_0[5|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|5]/row_en fgcell_amp_MiM_cap_1_10_0[6|4]/vsrc fgcell_amp_MiM_cap_1_10_0[7|0]/vdd
+ fgcell_amp_MiM_cap_1_10_0[7|0]/vinj fgcell_amp_MiM_cap_1_10_0[5|0]/row_en fgcell_amp_MiM_cap_1_10_0[6|7]/vdd
+ fgcell_amp_MiM_cap_1_10_0[8|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|6]/vtun fgcell_amp_MiM_cap_1_10_0[3|9]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[9|0]/row_en fgcell_amp_MiM_cap_1_10_0[2|8]/vinj fgcell_amp_MiM_cap_1_10_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|6]/row_en fgcell_amp_MiM_cap_1_10_0[6|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|5]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|0]/row_en fgcell_amp_MiM_cap_1_10_0[0|3]/vinj
+ fgcell_amp_MiM_cap_1_10_0[6|8]/row_en_b fgcell_amp_MiM_cap_1_10_0[6|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|0]/vtun fgcell_amp_MiM_cap_1_10_0[8|5]/vinj fgcell_amp_MiM_cap_1_10_0[1|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|2]/vtun fgcell_amp_MiM_cap_1_10_0[2|0]/vdd fgcell_amp_MiM_cap_1_10_0[7|2]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[7|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|7]/vtun fgcell_amp_MiM_cap_1_10_0[9|0]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[5|6]/row_en fgcell_amp_MiM_cap_1_10_0[5|0]/vdd fgcell_amp_MiM_cap_1_10_0[6|5]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[2|8]/vdd fgcell_amp_MiM_cap_1_10_0[6|9]/vdd fgcell_amp_MiM_cap_1_10_0[8|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|5]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|8]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|6]/vtun fgcell_amp_MiM_cap_1_10_0[1|8]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|1]/row_en fgcell_amp_MiM_cap_1_10_0[8|4]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[2|2]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|1]/vinj fgcell_amp_MiM_cap_1_10_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|4]/vinj fgcell_amp_MiM_cap_1_10_0[8|6]/vinj fgcell_amp_MiM_cap_1_10_0[0|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|3]/vtun fgcell_amp_MiM_cap_1_10_0[4|7]/row_en fgcell_amp_MiM_cap_1_10_0[9|1]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[1|9]/vdd fgcell_amp_MiM_cap_1_10_0[2|9]/vinj fgcell_amp_MiM_cap_1_10_0[2|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|8]/vtun fgcell_amp_MiM_cap_1_10_0[1|1]/vdd fgcell_amp_MiM_cap_1_10_0[8|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|6]/vsrc fgcell_amp_MiM_cap_1_10_0[9|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|5]/vdd fgcell_amp_MiM_cap_1_10_0[1|7]/row_en fgcell_amp_MiM_cap_1_10_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[4|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|0]/vinj fgcell_amp_MiM_cap_1_10_0[8|2]/row_en fgcell_amp_MiM_cap_1_10_0[0|5]/vinj
+ fgcell_amp_MiM_cap_1_10_0[8|0]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[0|2]/vtun fgcell_amp_MiM_cap_1_10_0[8|7]/vinj
+ fgcell_amp_MiM_cap_1_10_0[8|4]/vtun fgcell_amp_MiM_cap_1_10_0[1|0]/vsrc fgcell_amp_MiM_cap_1_10_0[7|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|2]/vsrc fgcell_amp_MiM_cap_1_10_0[6|9]/vinj fgcell_amp_MiM_cap_1_10_0[1|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|8]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|5]/vdd fgcell_amp_MiM_cap_1_10_0[6|7]/vsrc fgcell_amp_MiM_cap_1_10_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|3]/vdd fgcell_amp_MiM_cap_1_10_0[9|9]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|7]/vdd
+ fgcell_amp_MiM_cap_1_10_0[7|2]/vinj fgcell_amp_MiM_cap_1_10_0[4|8]/row_en fgcell_amp_MiM_cap_1_10_0[6|4]/vdd
+ fgcell_amp_MiM_cap_1_10_0[7|3]/row_en fgcell_amp_MiM_cap_1_10_0[5|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[3|1]/vinj fgcell_amp_MiM_cap_1_10_0[7|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|6]/vinj fgcell_amp_MiM_cap_1_10_0[8|8]/vinj fgcell_amp_MiM_cap_1_10_0[0|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|3]/vtun fgcell_amp_MiM_cap_1_10_0[8|5]/vtun fgcell_amp_MiM_cap_1_10_0[4|9]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|1]/vsrc fgcell_amp_MiM_cap_1_10_0[9|3]/vsrc fgcell_amp_MiM_cap_1_10_0[8|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[4|3]/row_en fgcell_amp_MiM_cap_1_10_0[8|0]/row_en_b fgcell_amp_MiM_cap_1_10_0[3|3]/vdd
+ fgcell_amp_MiM_cap_1_10_0[1|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|8]/vsrc fgcell_amp_MiM_cap_1_10_0[5|3]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[7|1]/vdd fgcell_amp_MiM_cap_1_10_0[3|9]/row_en fgcell_amp_MiM_cap_1_10_0[1|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|6]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|4]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[0|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[7|9]/row_en fgcell_amp_MiM_cap_1_10_0[3|0]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[2|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|2]/vinj fgcell_amp_MiM_cap_1_10_0[8|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|7]/vinj fgcell_amp_MiM_cap_1_10_0[0|3]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|4]/vtun fgcell_amp_MiM_cap_1_10_0[8|9]/vinj fgcell_amp_MiM_cap_1_10_0[3|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|6]/vtun fgcell_amp_MiM_cap_1_10_0[1|2]/vsrc fgcell_amp_MiM_cap_1_10_0[7|3]/vinj
+ fgcell_amp_MiM_cap_1_10_0[1|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|4]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[2|1]/vdd fgcell_amp_MiM_cap_1_10_0[7|4]/row_en fgcell_amp_MiM_cap_1_10_0[2|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|9]/vtun fgcell_amp_MiM_cap_1_10_0[6|9]/vsrc fgcell_amp_MiM_cap_1_10_0[4|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[8|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|4]/row_en fgcell_amp_MiM_cap_1_10_0[4|0]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|3]/vinj fgcell_amp_MiM_cap_1_10_0[3|0]/vtun fgcell_amp_MiM_cap_1_10_0[4|3]/vdd
+ fgcell_amp_MiM_cap_1_10_0[0|8]/vinj fgcell_amp_MiM_cap_1_10_0[0|5]/vtun fgcell_amp_MiM_cap_1_10_0[8|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|5]/row_en fgcell_amp_MiM_cap_1_10_0[4|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[1|3]/vsrc fgcell_amp_MiM_cap_1_10_0[9|5]/vsrc fgcell_amp_MiM_cap_1_10_0[7|8]/vdd
+ fgcell_amp_MiM_cap_1_10_0[3|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|9]/vtun fgcell_amp_MiM_cap_1_10_0[5|8]/vdd
+ fgcell_amp_MiM_cap_1_10_0[9|6]/vdd fgcell_amp_MiM_cap_1_10_0[3|5]/row_en fgcell_amp_MiM_cap_1_10_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|2]/vtun fgcell_amp_MiM_cap_1_10_0[7|4]/vinj fgcell_amp_MiM_cap_1_10_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|4]/vinj fgcell_amp_MiM_cap_1_10_0[1|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|4]/vdd fgcell_amp_MiM_cap_1_10_0[8|4]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|9]/vinj
+ fgcell_amp_MiM_cap_1_10_0[0|6]/vtun fgcell_amp_MiM_cap_1_10_0[6|1]/vdd fgcell_amp_MiM_cap_1_10_0[5|7]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[9|6]/row_en fgcell_amp_MiM_cap_1_10_0[8|8]/vtun fgcell_amp_MiM_cap_1_10_0[1|4]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[0|8]/vdd fgcell_amp_MiM_cap_1_10_0[3|0]/row_en fgcell_amp_MiM_cap_1_10_0[7|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[9|6]/vsrc fgcell_amp_MiM_cap_1_10_0[3|9]/vdd fgcell_amp_MiM_cap_1_10_0[4|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|6]/vdd fgcell_amp_MiM_cap_1_10_0[6|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|4]/vdd fgcell_amp_MiM_cap_1_10_0[3|4]/row_en_b fgcell_amp_MiM_cap_1_10_0[0|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[6|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|6]/row_en fgcell_amp_MiM_cap_1_10_0[6|0]/vinj
+ fgcell_amp_MiM_cap_1_10_0[0|7]/row_en_b fgcell_amp_MiM_cap_1_10_0[9|1]/row_en fgcell_amp_MiM_cap_1_10_0[7|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|5]/vinj fgcell_amp_MiM_cap_1_10_0[3|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|6]/vsrc fgcell_amp_MiM_cap_1_10_0[1|1]/row_en_b fgcell_amp_MiM_cap_1_10_0[4|0]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[2|1]/row_en fgcell_amp_MiM_cap_1_10_0[0|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[0|7]/vtun fgcell_amp_MiM_cap_1_10_0[8|9]/vtun fgcell_amp_MiM_cap_1_10_0[1|5]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[9|7]/vsrc fgcell_amp_MiM_cap_1_10_0[6|1]/row_en fgcell_amp_MiM_cap_1_10_0[9|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|4]/vdd fgcell_amp_MiM_cap_1_10_0[7|5]/vinj fgcell_amp_MiM_cap_1_10_0[0|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_10_0[5|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[5|7]/vdd fgcell_amp_MiM_cap_1_10_0[7|2]/vdd
+ fgcell_amp_MiM_cap_1_10_0[3|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[6|1]/vinj fgcell_amp_MiM_cap_1_10_0[9|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|3]/vtun fgcell_amp_MiM_cap_1_10_0[3|6]/vinj
+ fgcell_amp_MiM_cap_1_10_0[2|7]/row_en fgcell_amp_MiM_cap_1_10_0[4|1]/vsrc fgcell_amp_MiM_cap_1_10_0[4|6]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[0|8]/vtun fgcell_amp_MiM_cap_1_10_0[3|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[5|2]/row_en fgcell_amp_MiM_cap_1_10_0[1|6]/vsrc fgcell_amp_MiM_cap_1_10_0[9|8]/vsrc
+ fgcell_amp_MiM_cap_1_10_0[2|2]/vdd fgcell_amp_MiM_cap_1_10_0[4|0]/vdd fgcell_amp_MiM_cap_1_10_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|9]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[1|8]/vdd fgcell_amp_MiM_cap_1_10_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|0]/vdd fgcell_amp_MiM_cap_1_10_0[6|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_10_0[2|2]/row_en fgcell_amp_MiM_cap_1_10_0[5|5]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[7|5]/vdd
+ VSUBS fgcell_amp_MiM_cap_1_10_0[0|0]/vinj fgcell_amp_MiM_cap_1_10_0[6|2]/vinj fgcell_amp_MiM_cap_1_10_0[8|8]/row_en_b
+ fgcell_amp_MiM_cap_1_10_0[1|8]/row_en fgcell_amp_MiM_cap_1_10_0[4|1]/x1/x2/vb fgcell_amp_MiM_cap_1_10_0[3|7]/vinj
Xfgcell_amp_MiM_cap_1_10_0[0|0] fgcell_amp_MiM_cap_1_10_0[0|0]/vinj fgcell_amp_MiM_cap_1_10_0[0|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|0]/vdd fgcell_amp_MiM_cap_1_10_0[0|0]/vsrc fgcell_amp_MiM_cap_1_10_0[0|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|0] fgcell_amp_MiM_cap_1_10_0[1|0]/vinj fgcell_amp_MiM_cap_1_10_0[1|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|0]/vdd fgcell_amp_MiM_cap_1_10_0[1|0]/vsrc fgcell_amp_MiM_cap_1_10_0[1|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|0] fgcell_amp_MiM_cap_1_10_0[2|0]/vinj fgcell_amp_MiM_cap_1_10_0[2|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|0]/vdd fgcell_amp_MiM_cap_1_10_0[2|0]/vsrc fgcell_amp_MiM_cap_1_10_0[2|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|0] fgcell_amp_MiM_cap_1_10_0[3|0]/vinj fgcell_amp_MiM_cap_1_10_0[3|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|0]/vdd fgcell_amp_MiM_cap_1_10_0[3|0]/vsrc fgcell_amp_MiM_cap_1_10_0[3|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|0] fgcell_amp_MiM_cap_1_10_0[4|0]/vinj fgcell_amp_MiM_cap_1_10_0[4|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|0]/vdd fgcell_amp_MiM_cap_1_10_0[4|0]/vsrc fgcell_amp_MiM_cap_1_10_0[4|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|0] fgcell_amp_MiM_cap_1_10_0[5|0]/vinj fgcell_amp_MiM_cap_1_10_0[5|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|0]/vdd fgcell_amp_MiM_cap_1_10_0[5|0]/vsrc fgcell_amp_MiM_cap_1_10_0[5|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|0] fgcell_amp_MiM_cap_1_10_0[6|0]/vinj fgcell_amp_MiM_cap_1_10_0[6|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|0]/vdd fgcell_amp_MiM_cap_1_10_0[6|0]/vsrc fgcell_amp_MiM_cap_1_10_0[6|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|0] fgcell_amp_MiM_cap_1_10_0[7|0]/vinj fgcell_amp_MiM_cap_1_10_0[7|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|0]/vdd fgcell_amp_MiM_cap_1_10_0[7|0]/vsrc fgcell_amp_MiM_cap_1_10_0[7|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|0] fgcell_amp_MiM_cap_1_10_0[8|0]/vinj fgcell_amp_MiM_cap_1_10_0[8|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|0]/vdd fgcell_amp_MiM_cap_1_10_0[8|0]/vsrc fgcell_amp_MiM_cap_1_10_0[8|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|0] fgcell_amp_MiM_cap_1_10_0[9|0]/vinj fgcell_amp_MiM_cap_1_10_0[9|0]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|0]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|0]/vdd fgcell_amp_MiM_cap_1_10_0[9|0]/vsrc fgcell_amp_MiM_cap_1_10_0[9|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|1] fgcell_amp_MiM_cap_1_10_0[0|1]/vinj fgcell_amp_MiM_cap_1_10_0[0|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|1]/vdd fgcell_amp_MiM_cap_1_10_0[0|1]/vsrc fgcell_amp_MiM_cap_1_10_0[0|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|1] fgcell_amp_MiM_cap_1_10_0[1|1]/vinj fgcell_amp_MiM_cap_1_10_0[1|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|1]/vdd fgcell_amp_MiM_cap_1_10_0[1|1]/vsrc fgcell_amp_MiM_cap_1_10_0[1|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|1] fgcell_amp_MiM_cap_1_10_0[2|1]/vinj fgcell_amp_MiM_cap_1_10_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|1]/vdd fgcell_amp_MiM_cap_1_10_0[2|1]/vsrc fgcell_amp_MiM_cap_1_10_0[2|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|1] fgcell_amp_MiM_cap_1_10_0[3|1]/vinj fgcell_amp_MiM_cap_1_10_0[3|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|1]/vdd fgcell_amp_MiM_cap_1_10_0[3|1]/vsrc fgcell_amp_MiM_cap_1_10_0[3|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|1] fgcell_amp_MiM_cap_1_10_0[4|1]/vinj fgcell_amp_MiM_cap_1_10_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|1]/vdd fgcell_amp_MiM_cap_1_10_0[4|1]/vsrc fgcell_amp_MiM_cap_1_10_0[4|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|1] fgcell_amp_MiM_cap_1_10_0[5|1]/vinj fgcell_amp_MiM_cap_1_10_0[5|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|1]/vdd fgcell_amp_MiM_cap_1_10_0[5|1]/vsrc fgcell_amp_MiM_cap_1_10_0[5|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|1] fgcell_amp_MiM_cap_1_10_0[6|1]/vinj fgcell_amp_MiM_cap_1_10_0[6|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|1]/vdd fgcell_amp_MiM_cap_1_10_0[6|1]/vsrc fgcell_amp_MiM_cap_1_10_0[6|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|1] fgcell_amp_MiM_cap_1_10_0[7|1]/vinj fgcell_amp_MiM_cap_1_10_0[7|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|1]/vdd fgcell_amp_MiM_cap_1_10_0[7|1]/vsrc fgcell_amp_MiM_cap_1_10_0[7|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|1] fgcell_amp_MiM_cap_1_10_0[8|1]/vinj fgcell_amp_MiM_cap_1_10_0[8|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|1]/vdd fgcell_amp_MiM_cap_1_10_0[8|1]/vsrc fgcell_amp_MiM_cap_1_10_0[8|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|1] fgcell_amp_MiM_cap_1_10_0[9|1]/vinj fgcell_amp_MiM_cap_1_10_0[9|1]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|1]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|1]/vdd fgcell_amp_MiM_cap_1_10_0[9|1]/vsrc fgcell_amp_MiM_cap_1_10_0[9|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|2] fgcell_amp_MiM_cap_1_10_0[0|2]/vinj fgcell_amp_MiM_cap_1_10_0[0|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|2]/vdd fgcell_amp_MiM_cap_1_10_0[0|2]/vsrc fgcell_amp_MiM_cap_1_10_0[0|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|2] fgcell_amp_MiM_cap_1_10_0[1|2]/vinj fgcell_amp_MiM_cap_1_10_0[1|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|2]/vdd fgcell_amp_MiM_cap_1_10_0[1|2]/vsrc fgcell_amp_MiM_cap_1_10_0[1|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|2] fgcell_amp_MiM_cap_1_10_0[2|2]/vinj fgcell_amp_MiM_cap_1_10_0[2|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|2]/vdd fgcell_amp_MiM_cap_1_10_0[2|2]/vsrc fgcell_amp_MiM_cap_1_10_0[2|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|2] fgcell_amp_MiM_cap_1_10_0[3|2]/vinj fgcell_amp_MiM_cap_1_10_0[3|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|2]/vdd fgcell_amp_MiM_cap_1_10_0[3|2]/vsrc fgcell_amp_MiM_cap_1_10_0[3|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|2] fgcell_amp_MiM_cap_1_10_0[4|2]/vinj fgcell_amp_MiM_cap_1_10_0[4|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|2]/vdd fgcell_amp_MiM_cap_1_10_0[4|2]/vsrc fgcell_amp_MiM_cap_1_10_0[4|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|2] fgcell_amp_MiM_cap_1_10_0[5|2]/vinj fgcell_amp_MiM_cap_1_10_0[5|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|2]/vdd fgcell_amp_MiM_cap_1_10_0[5|2]/vsrc fgcell_amp_MiM_cap_1_10_0[5|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|2] fgcell_amp_MiM_cap_1_10_0[6|2]/vinj fgcell_amp_MiM_cap_1_10_0[6|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|2]/vdd fgcell_amp_MiM_cap_1_10_0[6|2]/vsrc fgcell_amp_MiM_cap_1_10_0[6|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|2] fgcell_amp_MiM_cap_1_10_0[7|2]/vinj fgcell_amp_MiM_cap_1_10_0[7|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|2]/vdd fgcell_amp_MiM_cap_1_10_0[7|2]/vsrc fgcell_amp_MiM_cap_1_10_0[7|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|2] fgcell_amp_MiM_cap_1_10_0[8|2]/vinj fgcell_amp_MiM_cap_1_10_0[8|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|2]/vdd fgcell_amp_MiM_cap_1_10_0[8|2]/vsrc fgcell_amp_MiM_cap_1_10_0[8|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|2] fgcell_amp_MiM_cap_1_10_0[9|2]/vinj fgcell_amp_MiM_cap_1_10_0[9|2]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|2]/vdd fgcell_amp_MiM_cap_1_10_0[9|2]/vsrc fgcell_amp_MiM_cap_1_10_0[9|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|3] fgcell_amp_MiM_cap_1_10_0[0|3]/vinj fgcell_amp_MiM_cap_1_10_0[0|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|3]/vdd fgcell_amp_MiM_cap_1_10_0[0|3]/vsrc fgcell_amp_MiM_cap_1_10_0[0|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|3] fgcell_amp_MiM_cap_1_10_0[1|3]/vinj fgcell_amp_MiM_cap_1_10_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|3]/vdd fgcell_amp_MiM_cap_1_10_0[1|3]/vsrc fgcell_amp_MiM_cap_1_10_0[1|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|3] fgcell_amp_MiM_cap_1_10_0[2|3]/vinj fgcell_amp_MiM_cap_1_10_0[2|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|3]/vdd fgcell_amp_MiM_cap_1_10_0[2|3]/vsrc fgcell_amp_MiM_cap_1_10_0[2|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|3] fgcell_amp_MiM_cap_1_10_0[3|3]/vinj fgcell_amp_MiM_cap_1_10_0[3|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|3]/vdd fgcell_amp_MiM_cap_1_10_0[3|3]/vsrc fgcell_amp_MiM_cap_1_10_0[3|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|3] fgcell_amp_MiM_cap_1_10_0[4|3]/vinj fgcell_amp_MiM_cap_1_10_0[4|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|3]/vdd fgcell_amp_MiM_cap_1_10_0[4|3]/vsrc fgcell_amp_MiM_cap_1_10_0[4|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|3] fgcell_amp_MiM_cap_1_10_0[5|3]/vinj fgcell_amp_MiM_cap_1_10_0[5|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|3]/vdd fgcell_amp_MiM_cap_1_10_0[5|3]/vsrc fgcell_amp_MiM_cap_1_10_0[5|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|3] fgcell_amp_MiM_cap_1_10_0[6|3]/vinj fgcell_amp_MiM_cap_1_10_0[6|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|3]/vdd fgcell_amp_MiM_cap_1_10_0[6|3]/vsrc fgcell_amp_MiM_cap_1_10_0[6|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|3] fgcell_amp_MiM_cap_1_10_0[7|3]/vinj fgcell_amp_MiM_cap_1_10_0[7|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|3]/vdd fgcell_amp_MiM_cap_1_10_0[7|3]/vsrc fgcell_amp_MiM_cap_1_10_0[7|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|3] fgcell_amp_MiM_cap_1_10_0[8|3]/vinj fgcell_amp_MiM_cap_1_10_0[8|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|3]/vdd fgcell_amp_MiM_cap_1_10_0[8|3]/vsrc fgcell_amp_MiM_cap_1_10_0[8|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|3] fgcell_amp_MiM_cap_1_10_0[9|3]/vinj fgcell_amp_MiM_cap_1_10_0[9|3]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|3]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|3]/vdd fgcell_amp_MiM_cap_1_10_0[9|3]/vsrc fgcell_amp_MiM_cap_1_10_0[9|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|4] fgcell_amp_MiM_cap_1_10_0[0|4]/vinj fgcell_amp_MiM_cap_1_10_0[0|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|4]/vdd fgcell_amp_MiM_cap_1_10_0[0|4]/vsrc fgcell_amp_MiM_cap_1_10_0[0|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|4] fgcell_amp_MiM_cap_1_10_0[1|4]/vinj fgcell_amp_MiM_cap_1_10_0[1|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|4]/vdd fgcell_amp_MiM_cap_1_10_0[1|4]/vsrc fgcell_amp_MiM_cap_1_10_0[1|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|4] fgcell_amp_MiM_cap_1_10_0[2|4]/vinj fgcell_amp_MiM_cap_1_10_0[2|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|4]/vdd fgcell_amp_MiM_cap_1_10_0[2|4]/vsrc fgcell_amp_MiM_cap_1_10_0[2|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|4] fgcell_amp_MiM_cap_1_10_0[3|4]/vinj fgcell_amp_MiM_cap_1_10_0[3|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|4]/vdd fgcell_amp_MiM_cap_1_10_0[3|4]/vsrc fgcell_amp_MiM_cap_1_10_0[3|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|4] fgcell_amp_MiM_cap_1_10_0[4|4]/vinj fgcell_amp_MiM_cap_1_10_0[4|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|4]/vdd fgcell_amp_MiM_cap_1_10_0[4|4]/vsrc fgcell_amp_MiM_cap_1_10_0[4|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|4] fgcell_amp_MiM_cap_1_10_0[5|4]/vinj fgcell_amp_MiM_cap_1_10_0[5|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|4]/vdd fgcell_amp_MiM_cap_1_10_0[5|4]/vsrc fgcell_amp_MiM_cap_1_10_0[5|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|4] fgcell_amp_MiM_cap_1_10_0[6|4]/vinj fgcell_amp_MiM_cap_1_10_0[6|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|4]/vdd fgcell_amp_MiM_cap_1_10_0[6|4]/vsrc fgcell_amp_MiM_cap_1_10_0[6|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|4] fgcell_amp_MiM_cap_1_10_0[7|4]/vinj fgcell_amp_MiM_cap_1_10_0[7|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|4]/vdd fgcell_amp_MiM_cap_1_10_0[7|4]/vsrc fgcell_amp_MiM_cap_1_10_0[7|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|4] fgcell_amp_MiM_cap_1_10_0[8|4]/vinj fgcell_amp_MiM_cap_1_10_0[8|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|4]/vdd fgcell_amp_MiM_cap_1_10_0[8|4]/vsrc fgcell_amp_MiM_cap_1_10_0[8|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|4] fgcell_amp_MiM_cap_1_10_0[9|4]/vinj fgcell_amp_MiM_cap_1_10_0[9|4]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|4]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|4]/vdd fgcell_amp_MiM_cap_1_10_0[9|4]/vsrc fgcell_amp_MiM_cap_1_10_0[9|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|5] fgcell_amp_MiM_cap_1_10_0[0|5]/vinj fgcell_amp_MiM_cap_1_10_0[0|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|5]/vdd fgcell_amp_MiM_cap_1_10_0[0|5]/vsrc fgcell_amp_MiM_cap_1_10_0[0|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|5] fgcell_amp_MiM_cap_1_10_0[1|5]/vinj fgcell_amp_MiM_cap_1_10_0[1|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|5]/vdd fgcell_amp_MiM_cap_1_10_0[1|5]/vsrc fgcell_amp_MiM_cap_1_10_0[1|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|5] fgcell_amp_MiM_cap_1_10_0[2|5]/vinj fgcell_amp_MiM_cap_1_10_0[2|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|5]/vdd fgcell_amp_MiM_cap_1_10_0[2|5]/vsrc fgcell_amp_MiM_cap_1_10_0[2|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|5] fgcell_amp_MiM_cap_1_10_0[3|5]/vinj fgcell_amp_MiM_cap_1_10_0[3|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|5]/vdd fgcell_amp_MiM_cap_1_10_0[3|5]/vsrc fgcell_amp_MiM_cap_1_10_0[3|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|5] fgcell_amp_MiM_cap_1_10_0[4|5]/vinj fgcell_amp_MiM_cap_1_10_0[4|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|5]/vdd fgcell_amp_MiM_cap_1_10_0[4|5]/vsrc fgcell_amp_MiM_cap_1_10_0[4|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|5] fgcell_amp_MiM_cap_1_10_0[5|5]/vinj fgcell_amp_MiM_cap_1_10_0[5|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|5]/vdd fgcell_amp_MiM_cap_1_10_0[5|5]/vsrc fgcell_amp_MiM_cap_1_10_0[5|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|5] fgcell_amp_MiM_cap_1_10_0[6|5]/vinj fgcell_amp_MiM_cap_1_10_0[6|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|5]/vdd fgcell_amp_MiM_cap_1_10_0[6|5]/vsrc fgcell_amp_MiM_cap_1_10_0[6|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|5] fgcell_amp_MiM_cap_1_10_0[7|5]/vinj fgcell_amp_MiM_cap_1_10_0[7|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|5]/vdd fgcell_amp_MiM_cap_1_10_0[7|5]/vsrc fgcell_amp_MiM_cap_1_10_0[7|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|5] fgcell_amp_MiM_cap_1_10_0[8|5]/vinj fgcell_amp_MiM_cap_1_10_0[8|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|5]/vdd fgcell_amp_MiM_cap_1_10_0[8|5]/vsrc fgcell_amp_MiM_cap_1_10_0[8|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|5] fgcell_amp_MiM_cap_1_10_0[9|5]/vinj fgcell_amp_MiM_cap_1_10_0[9|5]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|5]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|5]/vdd fgcell_amp_MiM_cap_1_10_0[9|5]/vsrc fgcell_amp_MiM_cap_1_10_0[9|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|6] fgcell_amp_MiM_cap_1_10_0[0|6]/vinj fgcell_amp_MiM_cap_1_10_0[0|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|6]/vdd fgcell_amp_MiM_cap_1_10_0[0|6]/vsrc fgcell_amp_MiM_cap_1_10_0[0|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|6] fgcell_amp_MiM_cap_1_10_0[1|6]/vinj fgcell_amp_MiM_cap_1_10_0[1|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|6]/vdd fgcell_amp_MiM_cap_1_10_0[1|6]/vsrc fgcell_amp_MiM_cap_1_10_0[1|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|6] fgcell_amp_MiM_cap_1_10_0[2|6]/vinj fgcell_amp_MiM_cap_1_10_0[2|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|6]/vdd fgcell_amp_MiM_cap_1_10_0[2|6]/vsrc fgcell_amp_MiM_cap_1_10_0[2|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|6] fgcell_amp_MiM_cap_1_10_0[3|6]/vinj fgcell_amp_MiM_cap_1_10_0[3|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|6]/vdd fgcell_amp_MiM_cap_1_10_0[3|6]/vsrc fgcell_amp_MiM_cap_1_10_0[3|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|6] fgcell_amp_MiM_cap_1_10_0[4|6]/vinj fgcell_amp_MiM_cap_1_10_0[4|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|6]/vdd fgcell_amp_MiM_cap_1_10_0[4|6]/vsrc fgcell_amp_MiM_cap_1_10_0[4|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|6] fgcell_amp_MiM_cap_1_10_0[5|6]/vinj fgcell_amp_MiM_cap_1_10_0[5|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|6]/vdd fgcell_amp_MiM_cap_1_10_0[5|6]/vsrc fgcell_amp_MiM_cap_1_10_0[5|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|6] fgcell_amp_MiM_cap_1_10_0[6|6]/vinj fgcell_amp_MiM_cap_1_10_0[6|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|6]/vdd fgcell_amp_MiM_cap_1_10_0[6|6]/vsrc fgcell_amp_MiM_cap_1_10_0[6|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|6] fgcell_amp_MiM_cap_1_10_0[7|6]/vinj fgcell_amp_MiM_cap_1_10_0[7|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|6]/vdd fgcell_amp_MiM_cap_1_10_0[7|6]/vsrc fgcell_amp_MiM_cap_1_10_0[7|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|6] fgcell_amp_MiM_cap_1_10_0[8|6]/vinj fgcell_amp_MiM_cap_1_10_0[8|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|6]/vdd fgcell_amp_MiM_cap_1_10_0[8|6]/vsrc fgcell_amp_MiM_cap_1_10_0[8|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|6] fgcell_amp_MiM_cap_1_10_0[9|6]/vinj fgcell_amp_MiM_cap_1_10_0[9|6]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|6]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|6]/vdd fgcell_amp_MiM_cap_1_10_0[9|6]/vsrc fgcell_amp_MiM_cap_1_10_0[9|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|7] fgcell_amp_MiM_cap_1_10_0[0|7]/vinj fgcell_amp_MiM_cap_1_10_0[0|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|7]/vdd fgcell_amp_MiM_cap_1_10_0[0|7]/vsrc fgcell_amp_MiM_cap_1_10_0[0|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|7] fgcell_amp_MiM_cap_1_10_0[1|7]/vinj fgcell_amp_MiM_cap_1_10_0[1|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|7]/vdd fgcell_amp_MiM_cap_1_10_0[1|7]/vsrc fgcell_amp_MiM_cap_1_10_0[1|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|7] fgcell_amp_MiM_cap_1_10_0[2|7]/vinj fgcell_amp_MiM_cap_1_10_0[2|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|7]/vdd fgcell_amp_MiM_cap_1_10_0[2|7]/vsrc fgcell_amp_MiM_cap_1_10_0[2|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|7] fgcell_amp_MiM_cap_1_10_0[3|7]/vinj fgcell_amp_MiM_cap_1_10_0[3|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|7]/vdd fgcell_amp_MiM_cap_1_10_0[3|7]/vsrc fgcell_amp_MiM_cap_1_10_0[3|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|7] fgcell_amp_MiM_cap_1_10_0[4|7]/vinj fgcell_amp_MiM_cap_1_10_0[4|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|7]/vdd fgcell_amp_MiM_cap_1_10_0[4|7]/vsrc fgcell_amp_MiM_cap_1_10_0[4|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|7] fgcell_amp_MiM_cap_1_10_0[5|7]/vinj fgcell_amp_MiM_cap_1_10_0[5|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|7]/vdd fgcell_amp_MiM_cap_1_10_0[5|7]/vsrc fgcell_amp_MiM_cap_1_10_0[5|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|7] fgcell_amp_MiM_cap_1_10_0[6|7]/vinj fgcell_amp_MiM_cap_1_10_0[6|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|7]/vdd fgcell_amp_MiM_cap_1_10_0[6|7]/vsrc fgcell_amp_MiM_cap_1_10_0[6|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|7] fgcell_amp_MiM_cap_1_10_0[7|7]/vinj fgcell_amp_MiM_cap_1_10_0[7|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|7]/vdd fgcell_amp_MiM_cap_1_10_0[7|7]/vsrc fgcell_amp_MiM_cap_1_10_0[7|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|7] fgcell_amp_MiM_cap_1_10_0[8|7]/vinj fgcell_amp_MiM_cap_1_10_0[8|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|7]/vdd fgcell_amp_MiM_cap_1_10_0[8|7]/vsrc fgcell_amp_MiM_cap_1_10_0[8|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|7] fgcell_amp_MiM_cap_1_10_0[9|7]/vinj fgcell_amp_MiM_cap_1_10_0[9|7]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|7]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|7]/vdd fgcell_amp_MiM_cap_1_10_0[9|7]/vsrc fgcell_amp_MiM_cap_1_10_0[9|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|8] fgcell_amp_MiM_cap_1_10_0[0|8]/vinj fgcell_amp_MiM_cap_1_10_0[0|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|8]/vdd fgcell_amp_MiM_cap_1_10_0[0|8]/vsrc fgcell_amp_MiM_cap_1_10_0[0|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|8] fgcell_amp_MiM_cap_1_10_0[1|8]/vinj fgcell_amp_MiM_cap_1_10_0[1|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|8]/vdd fgcell_amp_MiM_cap_1_10_0[1|8]/vsrc fgcell_amp_MiM_cap_1_10_0[1|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|8] fgcell_amp_MiM_cap_1_10_0[2|8]/vinj fgcell_amp_MiM_cap_1_10_0[2|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|8]/vdd fgcell_amp_MiM_cap_1_10_0[2|8]/vsrc fgcell_amp_MiM_cap_1_10_0[2|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|8] fgcell_amp_MiM_cap_1_10_0[3|8]/vinj fgcell_amp_MiM_cap_1_10_0[3|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|8]/vdd fgcell_amp_MiM_cap_1_10_0[3|8]/vsrc fgcell_amp_MiM_cap_1_10_0[3|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|8] fgcell_amp_MiM_cap_1_10_0[4|8]/vinj fgcell_amp_MiM_cap_1_10_0[4|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|8]/vdd fgcell_amp_MiM_cap_1_10_0[4|8]/vsrc fgcell_amp_MiM_cap_1_10_0[4|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|8] fgcell_amp_MiM_cap_1_10_0[5|8]/vinj fgcell_amp_MiM_cap_1_10_0[5|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|8]/vdd fgcell_amp_MiM_cap_1_10_0[5|8]/vsrc fgcell_amp_MiM_cap_1_10_0[5|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|8] fgcell_amp_MiM_cap_1_10_0[6|8]/vinj fgcell_amp_MiM_cap_1_10_0[6|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|8]/vdd fgcell_amp_MiM_cap_1_10_0[6|8]/vsrc fgcell_amp_MiM_cap_1_10_0[6|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|8] fgcell_amp_MiM_cap_1_10_0[7|8]/vinj fgcell_amp_MiM_cap_1_10_0[7|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|8]/vdd fgcell_amp_MiM_cap_1_10_0[7|8]/vsrc fgcell_amp_MiM_cap_1_10_0[7|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|8] fgcell_amp_MiM_cap_1_10_0[8|8]/vinj fgcell_amp_MiM_cap_1_10_0[8|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|8]/vdd fgcell_amp_MiM_cap_1_10_0[8|8]/vsrc fgcell_amp_MiM_cap_1_10_0[8|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|8] fgcell_amp_MiM_cap_1_10_0[9|8]/vinj fgcell_amp_MiM_cap_1_10_0[9|8]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|8]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|8]/vdd fgcell_amp_MiM_cap_1_10_0[9|8]/vsrc fgcell_amp_MiM_cap_1_10_0[9|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[0|9] fgcell_amp_MiM_cap_1_10_0[0|9]/vinj fgcell_amp_MiM_cap_1_10_0[0|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[0|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[0|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[0|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[0|9]/vdd fgcell_amp_MiM_cap_1_10_0[0|9]/vsrc fgcell_amp_MiM_cap_1_10_0[0|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[1|9] fgcell_amp_MiM_cap_1_10_0[1|9]/vinj fgcell_amp_MiM_cap_1_10_0[1|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[1|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[1|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[1|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[1|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[1|9]/vdd fgcell_amp_MiM_cap_1_10_0[1|9]/vsrc fgcell_amp_MiM_cap_1_10_0[1|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[2|9] fgcell_amp_MiM_cap_1_10_0[2|9]/vinj fgcell_amp_MiM_cap_1_10_0[2|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[2|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[2|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[2|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[2|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[2|9]/vdd fgcell_amp_MiM_cap_1_10_0[2|9]/vsrc fgcell_amp_MiM_cap_1_10_0[2|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[3|9] fgcell_amp_MiM_cap_1_10_0[3|9]/vinj fgcell_amp_MiM_cap_1_10_0[3|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[3|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[3|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[3|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[3|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[3|9]/vdd fgcell_amp_MiM_cap_1_10_0[3|9]/vsrc fgcell_amp_MiM_cap_1_10_0[3|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[4|9] fgcell_amp_MiM_cap_1_10_0[4|9]/vinj fgcell_amp_MiM_cap_1_10_0[4|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[4|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[4|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[4|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[4|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[4|9]/vdd fgcell_amp_MiM_cap_1_10_0[4|9]/vsrc fgcell_amp_MiM_cap_1_10_0[4|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[5|9] fgcell_amp_MiM_cap_1_10_0[5|9]/vinj fgcell_amp_MiM_cap_1_10_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[5|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[5|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[5|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[5|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[5|9]/vdd fgcell_amp_MiM_cap_1_10_0[5|9]/vsrc fgcell_amp_MiM_cap_1_10_0[5|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[6|9] fgcell_amp_MiM_cap_1_10_0[6|9]/vinj fgcell_amp_MiM_cap_1_10_0[6|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[6|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[6|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[6|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[6|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[6|9]/vdd fgcell_amp_MiM_cap_1_10_0[6|9]/vsrc fgcell_amp_MiM_cap_1_10_0[6|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[7|9] fgcell_amp_MiM_cap_1_10_0[7|9]/vinj fgcell_amp_MiM_cap_1_10_0[7|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[7|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[7|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[7|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[7|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[7|9]/vdd fgcell_amp_MiM_cap_1_10_0[7|9]/vsrc fgcell_amp_MiM_cap_1_10_0[7|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[8|9] fgcell_amp_MiM_cap_1_10_0[8|9]/vinj fgcell_amp_MiM_cap_1_10_0[8|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[8|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[8|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[8|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[8|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[8|9]/vdd fgcell_amp_MiM_cap_1_10_0[8|9]/vsrc fgcell_amp_MiM_cap_1_10_0[8|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
Xfgcell_amp_MiM_cap_1_10_0[9|9] fgcell_amp_MiM_cap_1_10_0[9|9]/vinj fgcell_amp_MiM_cap_1_10_0[9|9]/vtun
+ fgcell_amp_MiM_cap_1_10_0[9|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_10_0[9|9]/row_en
+ fgcell_amp_MiM_cap_1_10_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_10_0[9|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_10_0[9|9]/vdd fgcell_amp_MiM_cap_1_10_0[9|9]/vsrc fgcell_amp_MiM_cap_1_10_0[9|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_10
.ends

.subckt vb_divider VDD VGND vout_1v
X0 a_668_1320# a_556_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X1 a_332_1320# a_556_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X2 vout_1v a_1116_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X3 VGND a_444_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X4 a_892_1320# a_1116_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X5 a_892_1320# a_780_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X6 a_332_1320# a_220_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X7 vout_1v a_444_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X8 a_668_1320# a_780_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
X9 VDD a_220_220# VGND sky130_fd_pr__res_xhigh_po_0p35 l=3.5
.ends

.subckt fgcell_amp_MiM_cap_1_1 vinj vtun x1/tg5v0_0/vout row_en x1/x1/vctrl x1/x2/vb
+ vdd vsrc row_en_b VGND
Xx1 vtun x1/tg5v0_0/vout vdd x1/x2/v1 row_en vsrc x1/x1/vctrl row_en_b VGND vinj x1/x2/vb
+ fgcell_amp
X0 x1/x2/v1 VGND sky130_fd_pr__cap_mim_m3_1 l=1 w=1
.ends

.subckt array_core_block0 fgcell_amp_MiM_cap_1_1_0[0|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[6|0]/vtun fgcell_amp_MiM_cap_1_1_0[3|5]/vtun fgcell_amp_MiM_cap_1_1_0[5|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|3]/vsrc fgcell_amp_MiM_cap_1_1_0[8|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|8]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[1|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|0]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|8]/vinj
+ fgcell_amp_MiM_cap_1_1_0[6|4]/vinj fgcell_amp_MiM_cap_1_1_0[3|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|9]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[3|6]/vtun fgcell_amp_MiM_cap_1_1_0[4|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[4|4]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|3]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[1|9]/vsrc fgcell_amp_MiM_cap_1_1_0[1|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|5]/vinj fgcell_amp_MiM_cap_1_1_0[4|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[3|7]/vtun fgcell_amp_MiM_cap_1_1_0[7|0]/vsrc fgcell_amp_MiM_cap_1_1_0[9|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[4|5]/vsrc fgcell_amp_MiM_cap_1_1_0[2|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|9]/vinj fgcell_amp_MiM_cap_1_1_0[4|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|7]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|6]/vinj
+ fgcell_amp_MiM_cap_1_1_0[6|3]/vtun fgcell_amp_MiM_cap_1_1_0[7|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[7|1]/vsrc fgcell_amp_MiM_cap_1_1_0[3|8]/vtun fgcell_amp_MiM_cap_1_1_0[2|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|7]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[7|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[4|4]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|4]/vtun fgcell_amp_MiM_cap_1_1_0[3|4]/vdd
+ fgcell_amp_MiM_cap_1_1_0[6|7]/vinj fgcell_amp_MiM_cap_1_1_0[1|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|2]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[4|7]/vsrc fgcell_amp_MiM_cap_1_1_0[3|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|7]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[5|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|8]/vinj fgcell_amp_MiM_cap_1_1_0[3|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[6|5]/vtun fgcell_amp_MiM_cap_1_1_0[2|2]/vdd fgcell_amp_MiM_cap_1_1_0[7|3]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[0|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[6|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|8]/vsrc fgcell_amp_MiM_cap_1_1_0[3|9]/vtun fgcell_amp_MiM_cap_1_1_0[7|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[6|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|4]/vsrc fgcell_amp_MiM_cap_1_1_0[4|9]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[7|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|7]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[9|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[6|7]/vtun fgcell_amp_MiM_cap_1_1_0[2|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|5]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[2|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|2]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|1]/vtun fgcell_amp_MiM_cap_1_1_0[2|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|8]/vtun fgcell_amp_MiM_cap_1_1_0[1|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[3|5]/vdd fgcell_amp_MiM_cap_1_1_0[0|9]/vdd fgcell_amp_MiM_cap_1_1_0[7|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[5|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|3]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|0]/vsrc fgcell_amp_MiM_cap_1_1_0[5|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|3]/vdd fgcell_amp_MiM_cap_1_1_0[7|7]/vsrc fgcell_amp_MiM_cap_1_1_0[7|9]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[8|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|3]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|1]/vinj fgcell_amp_MiM_cap_1_1_0[8|4]/vdd
+ fgcell_amp_MiM_cap_1_1_0[1|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|1]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|0]/vinj
+ fgcell_amp_MiM_cap_1_1_0[3|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|8]/vsrc fgcell_amp_MiM_cap_1_1_0[1|0]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|2]/vinj
+ fgcell_amp_MiM_cap_1_1_0[4|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|4]/vtun fgcell_amp_MiM_cap_1_1_0[2|2]/vsrc fgcell_amp_MiM_cap_1_1_0[7|9]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[4|8]/vdd fgcell_amp_MiM_cap_1_1_0[4|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|3]/vinj fgcell_amp_MiM_cap_1_1_0[4|0]/vtun fgcell_amp_MiM_cap_1_1_0[1|1]/vinj
+ fgcell_amp_MiM_cap_1_1_0[1|4]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|5]/vtun fgcell_amp_MiM_cap_1_1_0[2|3]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[0|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[9|0]/vinj fgcell_amp_MiM_cap_1_1_0[9|8]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|6]/vdd fgcell_amp_MiM_cap_1_1_0[8|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|1]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[3|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|4]/vinj fgcell_amp_MiM_cap_1_1_0[6|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|4]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|4]/vsrc fgcell_amp_MiM_cap_1_1_0[1|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[5|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[4|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|4]/vdd fgcell_amp_MiM_cap_1_1_0[1|2]/vinj
+ fgcell_amp_MiM_cap_1_1_0[0|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[7|0]/vinj fgcell_amp_MiM_cap_1_1_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|5]/vinj fgcell_amp_MiM_cap_1_1_0[4|2]/vtun fgcell_amp_MiM_cap_1_1_0[3|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|0]/vsrc fgcell_amp_MiM_cap_1_1_0[9|1]/vinj fgcell_amp_MiM_cap_1_1_0[3|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|7]/vtun fgcell_amp_MiM_cap_1_1_0[2|5]/vsrc fgcell_amp_MiM_cap_1_1_0[2|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[3|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|1]/vinj fgcell_amp_MiM_cap_1_1_0[9|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[5|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|6]/vinj fgcell_amp_MiM_cap_1_1_0[6|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|3]/vtun fgcell_amp_MiM_cap_1_1_0[4|4]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|1]/vsrc fgcell_amp_MiM_cap_1_1_0[1|3]/vinj fgcell_amp_MiM_cap_1_1_0[3|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|0]/vdd fgcell_amp_MiM_cap_1_1_0[0|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[6|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|5]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|0]/vtun fgcell_amp_MiM_cap_1_1_0[6|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[9|2]/vinj fgcell_amp_MiM_cap_1_1_0[6|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[8|7]/vdd
+ fgcell_amp_MiM_cap_1_1_0[6|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|7]/vinj fgcell_amp_MiM_cap_1_1_0[7|2]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[4|4]/vtun fgcell_amp_MiM_cap_1_1_0[9|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|2]/vsrc fgcell_amp_MiM_cap_1_1_0[4|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|7]/vsrc fgcell_amp_MiM_cap_1_1_0[1|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|1]/vdd
+ fgcell_amp_MiM_cap_1_1_0[2|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|7]/vdd fgcell_amp_MiM_cap_1_1_0[2|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|4]/vinj
+ fgcell_amp_MiM_cap_1_1_0[7|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[7|0]/vtun fgcell_amp_MiM_cap_1_1_0[4|8]/vinj
+ fgcell_amp_MiM_cap_1_1_0[2|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|4]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[9|1]/vtun fgcell_amp_MiM_cap_1_1_0[5|3]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|3]/vinj fgcell_amp_MiM_cap_1_1_0[2|8]/vsrc fgcell_amp_MiM_cap_1_1_0[5|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[2|5]/vdd fgcell_amp_MiM_cap_1_1_0[6|3]/vdd fgcell_amp_MiM_cap_1_1_0[7|4]/vinj
+ fgcell_amp_MiM_cap_1_1_0[7|1]/vtun fgcell_amp_MiM_cap_1_1_0[8|8]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|9]/vinj
+ fgcell_amp_MiM_cap_1_1_0[7|4]/vdd fgcell_amp_MiM_cap_1_1_0[5|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|6]/vtun fgcell_amp_MiM_cap_1_1_0[5|4]/vsrc fgcell_amp_MiM_cap_1_1_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|9]/vsrc fgcell_amp_MiM_cap_1_1_0[1|5]/vinj
+ fgcell_amp_MiM_cap_1_1_0[9|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|0]/vdd fgcell_amp_MiM_cap_1_1_0[9|2]/vtun fgcell_amp_MiM_cap_1_1_0[7|6]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[7|5]/vinj fgcell_amp_MiM_cap_1_1_0[9|4]/vinj fgcell_amp_MiM_cap_1_1_0[9|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[8|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[4|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|0]/vsrc fgcell_amp_MiM_cap_1_1_0[8|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[8|4]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[5|5]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[2|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[7|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[8|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|6]/vinj fgcell_amp_MiM_cap_1_1_0[0|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|3]/vtun fgcell_amp_MiM_cap_1_1_0[8|1]/vsrc fgcell_amp_MiM_cap_1_1_0[1|6]/vinj
+ fgcell_amp_MiM_cap_1_1_0[1|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|6]/vsrc fgcell_amp_MiM_cap_1_1_0[7|1]/row_en fgcell_amp_MiM_cap_1_1_0[5|6]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|3]/vtun fgcell_amp_MiM_cap_1_1_0[4|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|8]/vdd fgcell_amp_MiM_cap_1_1_0[9|5]/vinj fgcell_amp_MiM_cap_1_1_0[0|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|8]/vdd fgcell_amp_MiM_cap_1_1_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|6]/vdd fgcell_amp_MiM_cap_1_1_0[7|7]/vinj fgcell_amp_MiM_cap_1_1_0[3|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|4]/vtun fgcell_amp_MiM_cap_1_1_0[0|0]/vsrc fgcell_amp_MiM_cap_1_1_0[4|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|9]/vtun fgcell_amp_MiM_cap_1_1_0[8|2]/vsrc fgcell_amp_MiM_cap_1_1_0[2|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|7]/vsrc fgcell_amp_MiM_cap_1_1_0[7|1]/vdd fgcell_amp_MiM_cap_1_1_0[4|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|2]/row_en fgcell_amp_MiM_cap_1_1_0[7|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[9|0]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|7]/vinj fgcell_amp_MiM_cap_1_1_0[2|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[1|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|0]/vinj fgcell_amp_MiM_cap_1_1_0[7|8]/vinj
+ fgcell_amp_MiM_cap_1_1_0[6|8]/row_en fgcell_amp_MiM_cap_1_1_0[7|5]/vtun fgcell_amp_MiM_cap_1_1_0[5|7]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|4]/vtun fgcell_amp_MiM_cap_1_1_0[0|1]/vsrc fgcell_amp_MiM_cap_1_1_0[8|3]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[7|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|6]/vinj fgcell_amp_MiM_cap_1_1_0[6|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|8]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[3|4]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[6|3]/row_en fgcell_amp_MiM_cap_1_1_0[0|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|4]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|1]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[2|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[5|2]/vdd fgcell_amp_MiM_cap_1_1_0[7|9]/vinj
+ fgcell_amp_MiM_cap_1_1_0[9|9]/row_en fgcell_amp_MiM_cap_1_1_0[7|6]/vtun fgcell_amp_MiM_cap_1_1_0[0|2]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[6|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[1|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|6]/vtun fgcell_amp_MiM_cap_1_1_0[8|4]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[1|8]/vinj fgcell_amp_MiM_cap_1_1_0[5|9]/vsrc fgcell_amp_MiM_cap_1_1_0[2|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|0]/vdd fgcell_amp_MiM_cap_1_1_0[2|1]/vinj fgcell_amp_MiM_cap_1_1_0[9|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|5]/vtun fgcell_amp_MiM_cap_1_1_0[0|2]/vdd fgcell_amp_MiM_cap_1_1_0[9|7]/vinj
+ fgcell_amp_MiM_cap_1_1_0[8|5]/vdd fgcell_amp_MiM_cap_1_1_0[6|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[6|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[3|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|4]/row_en fgcell_amp_MiM_cap_1_1_0[7|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|3]/vsrc fgcell_amp_MiM_cap_1_1_0[8|5]/vsrc fgcell_amp_MiM_cap_1_1_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|1]/vdd fgcell_amp_MiM_cap_1_1_0[8|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|1]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[3|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|9]/vinj fgcell_amp_MiM_cap_1_1_0[3|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[9|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[4|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[5|5]/row_en fgcell_amp_MiM_cap_1_1_0[7|7]/vdd fgcell_amp_MiM_cap_1_1_0[6|5]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[2|0]/vtun fgcell_amp_MiM_cap_1_1_0[7|8]/vtun fgcell_amp_MiM_cap_1_1_0[0|4]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[3|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|2]/vinj fgcell_amp_MiM_cap_1_1_0[3|8]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|6]/vtun fgcell_amp_MiM_cap_1_1_0[9|8]/vinj fgcell_amp_MiM_cap_1_1_0[4|2]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[2|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[5|0]/row_en fgcell_amp_MiM_cap_1_1_0[9|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|0]/vinj fgcell_amp_MiM_cap_1_1_0[1|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|7]/vdd
+ fgcell_amp_MiM_cap_1_1_0[4|6]/row_en fgcell_amp_MiM_cap_1_1_0[2|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|0]/vsrc fgcell_amp_MiM_cap_1_1_0[8|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|9]/vtun fgcell_amp_MiM_cap_1_1_0[6|4]/vdd fgcell_amp_MiM_cap_1_1_0[0|5]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|7]/vsrc fgcell_amp_MiM_cap_1_1_0[9|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|6]/row_en fgcell_amp_MiM_cap_1_1_0[4|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|1]/vinj fgcell_amp_MiM_cap_1_1_0[8|1]/row_en fgcell_amp_MiM_cap_1_1_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[7|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|3]/vinj fgcell_amp_MiM_cap_1_1_0[7|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|7]/vtun fgcell_amp_MiM_cap_1_1_0[5|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|1]/row_en fgcell_amp_MiM_cap_1_1_0[6|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|1]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|9]/vinj fgcell_amp_MiM_cap_1_1_0[5|3]/vdd fgcell_amp_MiM_cap_1_1_0[0|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[8|8]/vsrc fgcell_amp_MiM_cap_1_1_0[9|1]/vdd
+ fgcell_amp_MiM_cap_1_1_0[4|7]/row_en fgcell_amp_MiM_cap_1_1_0[7|2]/row_en fgcell_amp_MiM_cap_1_1_0[4|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|2]/vinj fgcell_amp_MiM_cap_1_1_0[0|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|2]/row_en fgcell_amp_MiM_cap_1_1_0[6|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|3]/vinj
+ fgcell_amp_MiM_cap_1_1_0[8|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|9]/vtun fgcell_amp_MiM_cap_1_1_0[3|2]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[4|1]/vdd fgcell_amp_MiM_cap_1_1_0[7|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|7]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|9]/vsrc fgcell_amp_MiM_cap_1_1_0[3|8]/row_en fgcell_amp_MiM_cap_1_1_0[1|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|4]/vinj fgcell_amp_MiM_cap_1_1_0[7|8]/row_en fgcell_amp_MiM_cap_1_1_0[1|9]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|8]/vtun fgcell_amp_MiM_cap_1_1_0[5|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|3]/vinj
+ fgcell_amp_MiM_cap_1_1_0[2|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|0]/vtun fgcell_amp_MiM_cap_1_1_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|3]/row_en fgcell_amp_MiM_cap_1_1_0[1|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|9]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/vsrc fgcell_amp_MiM_cap_1_1_0[7|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|8]/vsrc fgcell_amp_MiM_cap_1_1_0[7|8]/vdd
+ fgcell_amp_MiM_cap_1_1_0[7|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|3]/row_en fgcell_amp_MiM_cap_1_1_0[6|9]/row_en fgcell_amp_MiM_cap_1_1_0[6|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|1]/vdd fgcell_amp_MiM_cap_1_1_0[6|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|4]/vinj fgcell_amp_MiM_cap_1_1_0[3|9]/row_en fgcell_amp_MiM_cap_1_1_0[5|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|4]/row_en fgcell_amp_MiM_cap_1_1_0[2|3]/vtun fgcell_amp_MiM_cap_1_1_0[4|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|5]/vinj fgcell_amp_MiM_cap_1_1_0[2|8]/vdd fgcell_amp_MiM_cap_1_1_0[9|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|4]/vsrc fgcell_amp_MiM_cap_1_1_0[9|9]/vtun fgcell_amp_MiM_cap_1_1_0[6|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|9]/vsrc fgcell_amp_MiM_cap_1_1_0[8|5]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[7|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[3|4]/row_en fgcell_amp_MiM_cap_1_1_0[2|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|0]/vinj fgcell_amp_MiM_cap_1_1_0[0|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|5]/vinj fgcell_amp_MiM_cap_1_1_0[5|2]/vtun fgcell_amp_MiM_cap_1_1_0[7|7]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[9|5]/row_en fgcell_amp_MiM_cap_1_1_0[6|0]/vsrc fgcell_amp_MiM_cap_1_1_0[1|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[7|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|5]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[8|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|4]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|2]/vdd fgcell_amp_MiM_cap_1_1_0[2|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|0]/row_en fgcell_amp_MiM_cap_1_1_0[8|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[2|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|1]/vinj fgcell_amp_MiM_cap_1_1_0[2|6]/vinj fgcell_amp_MiM_cap_1_1_0[4|0]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|6]/vinj fgcell_amp_MiM_cap_1_1_0[5|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|0]/row_en fgcell_amp_MiM_cap_1_1_0[0|4]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|1]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[0|4]/vdd fgcell_amp_MiM_cap_1_1_0[7|5]/vdd fgcell_amp_MiM_cap_1_1_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|6]/vsrc fgcell_amp_MiM_cap_1_1_0[4|2]/vdd fgcell_amp_MiM_cap_1_1_0[5|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|6]/row_en fgcell_amp_MiM_cap_1_1_0[3|9]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|1]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[0|0]/vinj fgcell_amp_MiM_cap_1_1_0[8|2]/vinj
+ fgcell_amp_MiM_cap_1_1_0[0|1]/vdd fgcell_amp_MiM_cap_1_1_0[5|7]/vinj fgcell_amp_MiM_cap_1_1_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|4]/vtun fgcell_amp_MiM_cap_1_1_0[7|6]/vsrc fgcell_amp_MiM_cap_1_1_0[5|9]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[5|1]/row_en fgcell_amp_MiM_cap_1_1_0[6|2]/vsrc fgcell_amp_MiM_cap_1_1_0[3|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[9|1]/row_en fgcell_amp_MiM_cap_1_1_0[3|7]/vsrc fgcell_amp_MiM_cap_1_1_0[6|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[9|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|5]/vtun fgcell_amp_MiM_cap_1_1_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[2|7]/vinj fgcell_amp_MiM_cap_1_1_0[8|7]/row_en fgcell_amp_MiM_cap_1_1_0[6|6]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|1]/row_en fgcell_amp_MiM_cap_1_1_0[0|1]/vinj fgcell_amp_MiM_cap_1_1_0[8|3]/vinj
+ fgcell_amp_MiM_cap_1_1_0[1|7]/row_en fgcell_amp_MiM_cap_1_1_0[8|0]/vtun fgcell_amp_MiM_cap_1_1_0[5|8]/vinj
+ fgcell_amp_MiM_cap_1_1_0[8|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[5|5]/vtun fgcell_amp_MiM_cap_1_1_0[6|1]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|2]/row_en fgcell_amp_MiM_cap_1_1_0[6|3]/vsrc fgcell_amp_MiM_cap_1_1_0[0|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[3|8]/vsrc fgcell_amp_MiM_cap_1_1_0[2|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[5|4]/vdd fgcell_amp_MiM_cap_1_1_0[1|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|2]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[1|2]/row_en fgcell_amp_MiM_cap_1_1_0[6|7]/vdd fgcell_amp_MiM_cap_1_1_0[9|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|2]/row_en fgcell_amp_MiM_cap_1_1_0[3|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|9]/vdd fgcell_amp_MiM_cap_1_1_0[0|2]/vinj fgcell_amp_MiM_cap_1_1_0[8|4]/vinj
+ fgcell_amp_MiM_cap_1_1_0[4|8]/row_en fgcell_amp_MiM_cap_1_1_0[8|1]/vtun fgcell_amp_MiM_cap_1_1_0[2|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|6]/vtun fgcell_amp_MiM_cap_1_1_0[5|9]/vinj
+ fgcell_amp_MiM_cap_1_1_0[5|6]/vtun fgcell_amp_MiM_cap_1_1_0[2|8]/vinj fgcell_amp_MiM_cap_1_1_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|4]/vsrc fgcell_amp_MiM_cap_1_1_0[9|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[3|9]/vsrc fgcell_amp_MiM_cap_1_1_0[1|7]/vdd fgcell_amp_MiM_cap_1_1_0[1|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|5]/vdd fgcell_amp_MiM_cap_1_1_0[4|3]/row_en fgcell_amp_MiM_cap_1_1_0[5|5]/vdd
+ fgcell_amp_MiM_cap_1_1_0[2|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|2]/vdd
+ fgcell_amp_MiM_cap_1_1_0[8|3]/row_en fgcell_amp_MiM_cap_1_1_0[1|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[9|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|3]/vinj fgcell_amp_MiM_cap_1_1_0[0|0]/vtun fgcell_amp_MiM_cap_1_1_0[8|5]/vinj
+ fgcell_amp_MiM_cap_1_1_0[7|9]/row_en fgcell_amp_MiM_cap_1_1_0[8|2]/vtun fgcell_amp_MiM_cap_1_1_0[5|8]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|3]/row_en fgcell_amp_MiM_cap_1_1_0[6|6]/vtun fgcell_amp_MiM_cap_1_1_0[9|0]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[5|7]/vtun fgcell_amp_MiM_cap_1_1_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|5]/vsrc fgcell_amp_MiM_cap_1_1_0[0|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|9]/row_en fgcell_amp_MiM_cap_1_1_0[3|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[4|3]/vdd
+ fgcell_amp_MiM_cap_1_1_0[7|4]/row_en fgcell_amp_MiM_cap_1_1_0[2|7]/vtun fgcell_amp_MiM_cap_1_1_0[5|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[2|9]/vinj fgcell_amp_MiM_cap_1_1_0[8|1]/vdd fgcell_amp_MiM_cap_1_1_0[2|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|0]/vdd fgcell_amp_MiM_cap_1_1_0[0|4]/vinj fgcell_amp_MiM_cap_1_1_0[8|6]/vinj
+ fgcell_amp_MiM_cap_1_1_0[0|4]/row_en fgcell_amp_MiM_cap_1_1_0[8|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|3]/vtun fgcell_amp_MiM_cap_1_1_0[8|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[4|4]/row_en fgcell_amp_MiM_cap_1_1_0[5|8]/vtun fgcell_amp_MiM_cap_1_1_0[9|1]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|6]/vsrc fgcell_amp_MiM_cap_1_1_0[1|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[6|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[4|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|1]/vdd
+ fgcell_amp_MiM_cap_1_1_0[7|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[3|9]/row_en_b fgcell_amp_MiM_cap_1_1_0[8|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|3]/row_en_b fgcell_amp_MiM_cap_1_1_0[3|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|0]/vinj
+ fgcell_amp_MiM_cap_1_1_0[5|1]/vdd fgcell_amp_MiM_cap_1_1_0[6|9]/vinj fgcell_amp_MiM_cap_1_1_0[0|5]/vinj
+ fgcell_amp_MiM_cap_1_1_0[3|5]/row_en fgcell_amp_MiM_cap_1_1_0[0|2]/vtun fgcell_amp_MiM_cap_1_1_0[8|7]/vinj
+ fgcell_amp_MiM_cap_1_1_0[1|6]/row_en_b fgcell_amp_MiM_cap_1_1_0[1|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[8|4]/vtun fgcell_amp_MiM_cap_1_1_0[7|5]/row_en fgcell_amp_MiM_cap_1_1_0[1|0]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|2]/vsrc fgcell_amp_MiM_cap_1_1_0[7|2]/vinj fgcell_amp_MiM_cap_1_1_0[8|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[2|0]/row_en_b fgcell_amp_MiM_cap_1_1_0[2|8]/vtun fgcell_amp_MiM_cap_1_1_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|7]/vsrc fgcell_amp_MiM_cap_1_1_0[0|5]/row_en fgcell_amp_MiM_cap_1_1_0[3|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|8]/vdd fgcell_amp_MiM_cap_1_1_0[7|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|1]/vinj fgcell_amp_MiM_cap_1_1_0[1|2]/vdd
+ fgcell_amp_MiM_cap_1_1_0[0|6]/vinj fgcell_amp_MiM_cap_1_1_0[8|8]/vinj fgcell_amp_MiM_cap_1_1_0[6|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|3]/vtun fgcell_amp_MiM_cap_1_1_0[8|5]/vtun fgcell_amp_MiM_cap_1_1_0[0|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|7]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|5]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[1|1]/vsrc fgcell_amp_MiM_cap_1_1_0[9|3]/vsrc fgcell_amp_MiM_cap_1_1_0[4|7]/vdd
+ fgcell_amp_MiM_cap_1_1_0[6|8]/vsrc fgcell_amp_MiM_cap_1_1_0[1|8]/vdd fgcell_amp_MiM_cap_1_1_0[3|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[6|1]/row_en fgcell_amp_MiM_cap_1_1_0[4|0]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|6]/vdd fgcell_amp_MiM_cap_1_1_0[7|3]/vinj fgcell_amp_MiM_cap_1_1_0[5|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|2]/vinj fgcell_amp_MiM_cap_1_1_0[9|4]/vdd fgcell_amp_MiM_cap_1_1_0[2|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[5|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|0]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[2|9]/vtun fgcell_amp_MiM_cap_1_1_0[0|7]/vinj fgcell_amp_MiM_cap_1_1_0[9|7]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|4]/vtun fgcell_amp_MiM_cap_1_1_0[3|0]/vdd fgcell_amp_MiM_cap_1_1_0[8|9]/vinj
+ fgcell_amp_MiM_cap_1_1_0[7|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|6]/vtun fgcell_amp_MiM_cap_1_1_0[3|1]/row_en fgcell_amp_MiM_cap_1_1_0[1|2]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|4]/vsrc fgcell_amp_MiM_cap_1_1_0[0|8]/vdd fgcell_amp_MiM_cap_1_1_0[2|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|9]/vsrc fgcell_amp_MiM_cap_1_1_0[6|5]/vdd fgcell_amp_MiM_cap_1_1_0[7|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|6]/vdd
+ fgcell_amp_MiM_cap_1_1_0[6|7]/row_en fgcell_amp_MiM_cap_1_1_0[4|7]/row_en_b fgcell_amp_MiM_cap_1_1_0[7|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[6|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/vinj
+ fgcell_amp_MiM_cap_1_1_0[8|2]/vdd fgcell_amp_MiM_cap_1_1_0[3|0]/vtun fgcell_amp_MiM_cap_1_1_0[2|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|9]/vtun fgcell_amp_MiM_cap_1_1_0[0|8]/vinj fgcell_amp_MiM_cap_1_1_0[2|4]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[0|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|7]/vtun fgcell_amp_MiM_cap_1_1_0[6|2]/row_en fgcell_amp_MiM_cap_1_1_0[1|3]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[7|2]/vtun fgcell_amp_MiM_cap_1_1_0[9|5]/vsrc fgcell_amp_MiM_cap_1_1_0[5|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|1]/row_en_b fgcell_amp_MiM_cap_1_1_0[3|7]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[9|8]/row_en fgcell_amp_MiM_cap_1_1_0[8|6]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|2]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|4]/vinj fgcell_amp_MiM_cap_1_1_0[7|0]/vdd fgcell_amp_MiM_cap_1_1_0[9|6]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[7|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|1]/vtun fgcell_amp_MiM_cap_1_1_0[2|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[6|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|9]/vinj fgcell_amp_MiM_cap_1_1_0[3|2]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|3]/row_en fgcell_amp_MiM_cap_1_1_0[0|6]/vtun fgcell_amp_MiM_cap_1_1_0[8|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|4]/vsrc fgcell_amp_MiM_cap_1_1_0[9|3]/row_en fgcell_amp_MiM_cap_1_1_0[9|6]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[6|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|3]/row_en fgcell_amp_MiM_cap_1_1_0[0|6]/vsrc fgcell_amp_MiM_cap_1_1_0[2|0]/vdd
+ fgcell_amp_MiM_cap_1_1_0[4|4]/vdd fgcell_amp_MiM_cap_1_1_0[9|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|0]/vinj fgcell_amp_MiM_cap_1_1_0[1|9]/row_en fgcell_amp_MiM_cap_1_1_0[0|4]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|2]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|5]/vinj fgcell_amp_MiM_cap_1_1_0[6|9]/vdd
+ fgcell_amp_MiM_cap_1_1_0[7|9]/vdd fgcell_amp_MiM_cap_1_1_0[3|2]/vtun fgcell_amp_MiM_cap_1_1_0[5|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|0]/vsrc fgcell_amp_MiM_cap_1_1_0[8|4]/row_en fgcell_amp_MiM_cap_1_1_0[6|3]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|7]/vtun fgcell_amp_MiM_cap_1_1_0[8|9]/vtun fgcell_amp_MiM_cap_1_1_0[7|8]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[1|5]/vsrc fgcell_amp_MiM_cap_1_1_0[9|7]/vsrc fgcell_amp_MiM_cap_1_1_0[1|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[9|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[5|4]/row_en fgcell_amp_MiM_cap_1_1_0[0|5]/vdd fgcell_amp_MiM_cap_1_1_0[5|5]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[4|6]/vsrc fgcell_amp_MiM_cap_1_1_0[1|9]/vdd fgcell_amp_MiM_cap_1_1_0[6|1]/vinj
+ fgcell_amp_MiM_cap_1_1_0[6|2]/vdd fgcell_amp_MiM_cap_1_1_0[2|8]/row_en_b fgcell_amp_MiM_cap_1_1_0[3|6]/vinj
+ fgcell_amp_MiM_cap_1_1_0[5|7]/vdd fgcell_amp_MiM_cap_1_1_0[2|9]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[9|2]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[3|3]/vtun fgcell_amp_MiM_cap_1_1_0[9|5]/vdd
+ fgcell_amp_MiM_cap_1_1_0[3|2]/row_en_b fgcell_amp_MiM_cap_1_1_0[0|8]/vtun fgcell_amp_MiM_cap_1_1_0[4|1]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[9|7]/vdd fgcell_amp_MiM_cap_1_1_0[9|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[1|6]/vsrc fgcell_amp_MiM_cap_1_1_0[0|5]/row_en_b fgcell_amp_MiM_cap_1_1_0[9|8]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[4|5]/row_en fgcell_amp_MiM_cap_1_1_0[2|4]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[0|7]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[8|5]/row_en fgcell_amp_MiM_cap_1_1_0[0|7]/vdd
+ fgcell_amp_MiM_cap_1_1_0[5|7]/row_en fgcell_amp_MiM_cap_1_1_0[4|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|8]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[8|6]/vsrc fgcell_amp_MiM_cap_1_1_0[6|2]/vinj fgcell_amp_MiM_cap_1_1_0[4|5]/vdd
+ fgcell_amp_MiM_cap_1_1_0[8|0]/vdd fgcell_amp_MiM_cap_1_1_0[1|5]/row_en fgcell_amp_MiM_cap_1_1_0[3|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|3]/vdd fgcell_amp_MiM_cap_1_1_0[4|0]/row_en fgcell_amp_MiM_cap_1_1_0[4|2]/vsrc
+ fgcell_amp_MiM_cap_1_1_0[5|8]/vdd fgcell_amp_MiM_cap_1_1_0[0|9]/vtun fgcell_amp_MiM_cap_1_1_0[3|7]/vinj
+ fgcell_amp_MiM_cap_1_1_0[8|0]/row_en fgcell_amp_MiM_cap_1_1_0[1|7]/vsrc fgcell_amp_MiM_cap_1_1_0[9|9]/vsrc
+ VSUBS fgcell_amp_MiM_cap_1_1_0[4|0]/vinj fgcell_amp_MiM_cap_1_1_0[5|6]/row_en_b
+ fgcell_amp_MiM_cap_1_1_0[7|6]/row_en fgcell_amp_MiM_cap_1_1_0[5|5]/x1/tg5v0_0/vout
+ fgcell_amp_MiM_cap_1_1_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|3]/x1/x1/vctrl
+ fgcell_amp_MiM_cap_1_1_0[1|7]/x1/x2/vb fgcell_amp_MiM_cap_1_1_0[1|0]/row_en fgcell_amp_MiM_cap_1_1_0[1|5]/x1/x1/vctrl
Xfgcell_amp_MiM_cap_1_1_0[0|0] fgcell_amp_MiM_cap_1_1_0[0|0]/vinj fgcell_amp_MiM_cap_1_1_0[0|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|0]/vdd fgcell_amp_MiM_cap_1_1_0[0|0]/vsrc fgcell_amp_MiM_cap_1_1_0[0|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|0] fgcell_amp_MiM_cap_1_1_0[1|0]/vinj fgcell_amp_MiM_cap_1_1_0[1|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|0]/vdd fgcell_amp_MiM_cap_1_1_0[1|0]/vsrc fgcell_amp_MiM_cap_1_1_0[1|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|0] fgcell_amp_MiM_cap_1_1_0[2|0]/vinj fgcell_amp_MiM_cap_1_1_0[2|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|0]/vdd fgcell_amp_MiM_cap_1_1_0[2|0]/vsrc fgcell_amp_MiM_cap_1_1_0[2|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|0] fgcell_amp_MiM_cap_1_1_0[3|0]/vinj fgcell_amp_MiM_cap_1_1_0[3|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|0]/vdd fgcell_amp_MiM_cap_1_1_0[3|0]/vsrc fgcell_amp_MiM_cap_1_1_0[3|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|0] fgcell_amp_MiM_cap_1_1_0[4|0]/vinj fgcell_amp_MiM_cap_1_1_0[4|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|0]/vdd fgcell_amp_MiM_cap_1_1_0[4|0]/vsrc fgcell_amp_MiM_cap_1_1_0[4|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|0] fgcell_amp_MiM_cap_1_1_0[5|0]/vinj fgcell_amp_MiM_cap_1_1_0[5|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|0]/vdd fgcell_amp_MiM_cap_1_1_0[5|0]/vsrc fgcell_amp_MiM_cap_1_1_0[5|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|0] fgcell_amp_MiM_cap_1_1_0[6|0]/vinj fgcell_amp_MiM_cap_1_1_0[6|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|0]/vdd fgcell_amp_MiM_cap_1_1_0[6|0]/vsrc fgcell_amp_MiM_cap_1_1_0[6|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|0] fgcell_amp_MiM_cap_1_1_0[7|0]/vinj fgcell_amp_MiM_cap_1_1_0[7|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|0]/vdd fgcell_amp_MiM_cap_1_1_0[7|0]/vsrc fgcell_amp_MiM_cap_1_1_0[7|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|0] fgcell_amp_MiM_cap_1_1_0[8|0]/vinj fgcell_amp_MiM_cap_1_1_0[8|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|0]/vdd fgcell_amp_MiM_cap_1_1_0[8|0]/vsrc fgcell_amp_MiM_cap_1_1_0[8|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|0] fgcell_amp_MiM_cap_1_1_0[9|0]/vinj fgcell_amp_MiM_cap_1_1_0[9|0]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|0]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|0]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|0]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|0]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|0]/vdd fgcell_amp_MiM_cap_1_1_0[9|0]/vsrc fgcell_amp_MiM_cap_1_1_0[9|0]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|1] fgcell_amp_MiM_cap_1_1_0[0|1]/vinj fgcell_amp_MiM_cap_1_1_0[0|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|1]/vdd fgcell_amp_MiM_cap_1_1_0[0|1]/vsrc fgcell_amp_MiM_cap_1_1_0[0|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|1] fgcell_amp_MiM_cap_1_1_0[1|1]/vinj fgcell_amp_MiM_cap_1_1_0[1|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|1]/vdd fgcell_amp_MiM_cap_1_1_0[1|1]/vsrc fgcell_amp_MiM_cap_1_1_0[1|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|1] fgcell_amp_MiM_cap_1_1_0[2|1]/vinj fgcell_amp_MiM_cap_1_1_0[2|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|1]/vdd fgcell_amp_MiM_cap_1_1_0[2|1]/vsrc fgcell_amp_MiM_cap_1_1_0[2|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|1] fgcell_amp_MiM_cap_1_1_0[3|1]/vinj fgcell_amp_MiM_cap_1_1_0[3|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|1]/vdd fgcell_amp_MiM_cap_1_1_0[3|1]/vsrc fgcell_amp_MiM_cap_1_1_0[3|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|1] fgcell_amp_MiM_cap_1_1_0[4|1]/vinj fgcell_amp_MiM_cap_1_1_0[4|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|1]/vdd fgcell_amp_MiM_cap_1_1_0[4|1]/vsrc fgcell_amp_MiM_cap_1_1_0[4|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|1] fgcell_amp_MiM_cap_1_1_0[5|1]/vinj fgcell_amp_MiM_cap_1_1_0[5|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|1]/vdd fgcell_amp_MiM_cap_1_1_0[5|1]/vsrc fgcell_amp_MiM_cap_1_1_0[5|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|1] fgcell_amp_MiM_cap_1_1_0[6|1]/vinj fgcell_amp_MiM_cap_1_1_0[6|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|1]/vdd fgcell_amp_MiM_cap_1_1_0[6|1]/vsrc fgcell_amp_MiM_cap_1_1_0[6|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|1] fgcell_amp_MiM_cap_1_1_0[7|1]/vinj fgcell_amp_MiM_cap_1_1_0[7|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|1]/vdd fgcell_amp_MiM_cap_1_1_0[7|1]/vsrc fgcell_amp_MiM_cap_1_1_0[7|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|1] fgcell_amp_MiM_cap_1_1_0[8|1]/vinj fgcell_amp_MiM_cap_1_1_0[8|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|1]/vdd fgcell_amp_MiM_cap_1_1_0[8|1]/vsrc fgcell_amp_MiM_cap_1_1_0[8|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|1] fgcell_amp_MiM_cap_1_1_0[9|1]/vinj fgcell_amp_MiM_cap_1_1_0[9|1]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|1]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|1]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|1]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|1]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|1]/vdd fgcell_amp_MiM_cap_1_1_0[9|1]/vsrc fgcell_amp_MiM_cap_1_1_0[9|1]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|2] fgcell_amp_MiM_cap_1_1_0[0|2]/vinj fgcell_amp_MiM_cap_1_1_0[0|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|2]/vdd fgcell_amp_MiM_cap_1_1_0[0|2]/vsrc fgcell_amp_MiM_cap_1_1_0[0|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|2] fgcell_amp_MiM_cap_1_1_0[1|2]/vinj fgcell_amp_MiM_cap_1_1_0[1|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|2]/vdd fgcell_amp_MiM_cap_1_1_0[1|2]/vsrc fgcell_amp_MiM_cap_1_1_0[1|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|2] fgcell_amp_MiM_cap_1_1_0[2|2]/vinj fgcell_amp_MiM_cap_1_1_0[2|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|2]/vdd fgcell_amp_MiM_cap_1_1_0[2|2]/vsrc fgcell_amp_MiM_cap_1_1_0[2|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|2] fgcell_amp_MiM_cap_1_1_0[3|2]/vinj fgcell_amp_MiM_cap_1_1_0[3|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|2]/vdd fgcell_amp_MiM_cap_1_1_0[3|2]/vsrc fgcell_amp_MiM_cap_1_1_0[3|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|2] fgcell_amp_MiM_cap_1_1_0[4|2]/vinj fgcell_amp_MiM_cap_1_1_0[4|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|2]/vdd fgcell_amp_MiM_cap_1_1_0[4|2]/vsrc fgcell_amp_MiM_cap_1_1_0[4|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|2] fgcell_amp_MiM_cap_1_1_0[5|2]/vinj fgcell_amp_MiM_cap_1_1_0[5|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|2]/vdd fgcell_amp_MiM_cap_1_1_0[5|2]/vsrc fgcell_amp_MiM_cap_1_1_0[5|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|2] fgcell_amp_MiM_cap_1_1_0[6|2]/vinj fgcell_amp_MiM_cap_1_1_0[6|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|2]/vdd fgcell_amp_MiM_cap_1_1_0[6|2]/vsrc fgcell_amp_MiM_cap_1_1_0[6|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|2] fgcell_amp_MiM_cap_1_1_0[7|2]/vinj fgcell_amp_MiM_cap_1_1_0[7|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|2]/vdd fgcell_amp_MiM_cap_1_1_0[7|2]/vsrc fgcell_amp_MiM_cap_1_1_0[7|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|2] fgcell_amp_MiM_cap_1_1_0[8|2]/vinj fgcell_amp_MiM_cap_1_1_0[8|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|2]/vdd fgcell_amp_MiM_cap_1_1_0[8|2]/vsrc fgcell_amp_MiM_cap_1_1_0[8|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|2] fgcell_amp_MiM_cap_1_1_0[9|2]/vinj fgcell_amp_MiM_cap_1_1_0[9|2]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|2]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|2]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|2]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|2]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|2]/vdd fgcell_amp_MiM_cap_1_1_0[9|2]/vsrc fgcell_amp_MiM_cap_1_1_0[9|2]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|3] fgcell_amp_MiM_cap_1_1_0[0|3]/vinj fgcell_amp_MiM_cap_1_1_0[0|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|3]/vdd fgcell_amp_MiM_cap_1_1_0[0|3]/vsrc fgcell_amp_MiM_cap_1_1_0[0|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|3] fgcell_amp_MiM_cap_1_1_0[1|3]/vinj fgcell_amp_MiM_cap_1_1_0[1|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|3]/vdd fgcell_amp_MiM_cap_1_1_0[1|3]/vsrc fgcell_amp_MiM_cap_1_1_0[1|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|3] fgcell_amp_MiM_cap_1_1_0[2|3]/vinj fgcell_amp_MiM_cap_1_1_0[2|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|3]/vdd fgcell_amp_MiM_cap_1_1_0[2|3]/vsrc fgcell_amp_MiM_cap_1_1_0[2|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|3] fgcell_amp_MiM_cap_1_1_0[3|3]/vinj fgcell_amp_MiM_cap_1_1_0[3|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|3]/vdd fgcell_amp_MiM_cap_1_1_0[3|3]/vsrc fgcell_amp_MiM_cap_1_1_0[3|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|3] fgcell_amp_MiM_cap_1_1_0[4|3]/vinj fgcell_amp_MiM_cap_1_1_0[4|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|3]/vdd fgcell_amp_MiM_cap_1_1_0[4|3]/vsrc fgcell_amp_MiM_cap_1_1_0[4|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|3] fgcell_amp_MiM_cap_1_1_0[5|3]/vinj fgcell_amp_MiM_cap_1_1_0[5|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|3]/vdd fgcell_amp_MiM_cap_1_1_0[5|3]/vsrc fgcell_amp_MiM_cap_1_1_0[5|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|3] fgcell_amp_MiM_cap_1_1_0[6|3]/vinj fgcell_amp_MiM_cap_1_1_0[6|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|3]/vdd fgcell_amp_MiM_cap_1_1_0[6|3]/vsrc fgcell_amp_MiM_cap_1_1_0[6|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|3] fgcell_amp_MiM_cap_1_1_0[7|3]/vinj fgcell_amp_MiM_cap_1_1_0[7|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|3]/vdd fgcell_amp_MiM_cap_1_1_0[7|3]/vsrc fgcell_amp_MiM_cap_1_1_0[7|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|3] fgcell_amp_MiM_cap_1_1_0[8|3]/vinj fgcell_amp_MiM_cap_1_1_0[8|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|3]/vdd fgcell_amp_MiM_cap_1_1_0[8|3]/vsrc fgcell_amp_MiM_cap_1_1_0[8|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|3] fgcell_amp_MiM_cap_1_1_0[9|3]/vinj fgcell_amp_MiM_cap_1_1_0[9|3]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|3]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|3]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|3]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|3]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|3]/vdd fgcell_amp_MiM_cap_1_1_0[9|3]/vsrc fgcell_amp_MiM_cap_1_1_0[9|3]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|4] fgcell_amp_MiM_cap_1_1_0[0|4]/vinj fgcell_amp_MiM_cap_1_1_0[0|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|4]/vdd fgcell_amp_MiM_cap_1_1_0[0|4]/vsrc fgcell_amp_MiM_cap_1_1_0[0|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|4] fgcell_amp_MiM_cap_1_1_0[1|4]/vinj fgcell_amp_MiM_cap_1_1_0[1|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|4]/vdd fgcell_amp_MiM_cap_1_1_0[1|4]/vsrc fgcell_amp_MiM_cap_1_1_0[1|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|4] fgcell_amp_MiM_cap_1_1_0[2|4]/vinj fgcell_amp_MiM_cap_1_1_0[2|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|4]/vdd fgcell_amp_MiM_cap_1_1_0[2|4]/vsrc fgcell_amp_MiM_cap_1_1_0[2|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|4] fgcell_amp_MiM_cap_1_1_0[3|4]/vinj fgcell_amp_MiM_cap_1_1_0[3|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|4]/vdd fgcell_amp_MiM_cap_1_1_0[3|4]/vsrc fgcell_amp_MiM_cap_1_1_0[3|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|4] fgcell_amp_MiM_cap_1_1_0[4|4]/vinj fgcell_amp_MiM_cap_1_1_0[4|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|4]/vdd fgcell_amp_MiM_cap_1_1_0[4|4]/vsrc fgcell_amp_MiM_cap_1_1_0[4|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|4] fgcell_amp_MiM_cap_1_1_0[5|4]/vinj fgcell_amp_MiM_cap_1_1_0[5|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|4]/vdd fgcell_amp_MiM_cap_1_1_0[5|4]/vsrc fgcell_amp_MiM_cap_1_1_0[5|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|4] fgcell_amp_MiM_cap_1_1_0[6|4]/vinj fgcell_amp_MiM_cap_1_1_0[6|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|4]/vdd fgcell_amp_MiM_cap_1_1_0[6|4]/vsrc fgcell_amp_MiM_cap_1_1_0[6|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|4] fgcell_amp_MiM_cap_1_1_0[7|4]/vinj fgcell_amp_MiM_cap_1_1_0[7|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|4]/vdd fgcell_amp_MiM_cap_1_1_0[7|4]/vsrc fgcell_amp_MiM_cap_1_1_0[7|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|4] fgcell_amp_MiM_cap_1_1_0[8|4]/vinj fgcell_amp_MiM_cap_1_1_0[8|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|4]/vdd fgcell_amp_MiM_cap_1_1_0[8|4]/vsrc fgcell_amp_MiM_cap_1_1_0[8|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|4] fgcell_amp_MiM_cap_1_1_0[9|4]/vinj fgcell_amp_MiM_cap_1_1_0[9|4]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|4]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|4]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|4]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|4]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|4]/vdd fgcell_amp_MiM_cap_1_1_0[9|4]/vsrc fgcell_amp_MiM_cap_1_1_0[9|4]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|5] fgcell_amp_MiM_cap_1_1_0[0|5]/vinj fgcell_amp_MiM_cap_1_1_0[0|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|5]/vdd fgcell_amp_MiM_cap_1_1_0[0|5]/vsrc fgcell_amp_MiM_cap_1_1_0[0|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|5] fgcell_amp_MiM_cap_1_1_0[1|5]/vinj fgcell_amp_MiM_cap_1_1_0[1|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|5]/vdd fgcell_amp_MiM_cap_1_1_0[1|5]/vsrc fgcell_amp_MiM_cap_1_1_0[1|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|5] fgcell_amp_MiM_cap_1_1_0[2|5]/vinj fgcell_amp_MiM_cap_1_1_0[2|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|5]/vdd fgcell_amp_MiM_cap_1_1_0[2|5]/vsrc fgcell_amp_MiM_cap_1_1_0[2|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|5] fgcell_amp_MiM_cap_1_1_0[3|5]/vinj fgcell_amp_MiM_cap_1_1_0[3|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|5]/vdd fgcell_amp_MiM_cap_1_1_0[3|5]/vsrc fgcell_amp_MiM_cap_1_1_0[3|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|5] fgcell_amp_MiM_cap_1_1_0[4|5]/vinj fgcell_amp_MiM_cap_1_1_0[4|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|5]/vdd fgcell_amp_MiM_cap_1_1_0[4|5]/vsrc fgcell_amp_MiM_cap_1_1_0[4|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|5] fgcell_amp_MiM_cap_1_1_0[5|5]/vinj fgcell_amp_MiM_cap_1_1_0[5|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|5]/vdd fgcell_amp_MiM_cap_1_1_0[5|5]/vsrc fgcell_amp_MiM_cap_1_1_0[5|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|5] fgcell_amp_MiM_cap_1_1_0[6|5]/vinj fgcell_amp_MiM_cap_1_1_0[6|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|5]/vdd fgcell_amp_MiM_cap_1_1_0[6|5]/vsrc fgcell_amp_MiM_cap_1_1_0[6|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|5] fgcell_amp_MiM_cap_1_1_0[7|5]/vinj fgcell_amp_MiM_cap_1_1_0[7|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|5]/vdd fgcell_amp_MiM_cap_1_1_0[7|5]/vsrc fgcell_amp_MiM_cap_1_1_0[7|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|5] fgcell_amp_MiM_cap_1_1_0[8|5]/vinj fgcell_amp_MiM_cap_1_1_0[8|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|5]/vdd fgcell_amp_MiM_cap_1_1_0[8|5]/vsrc fgcell_amp_MiM_cap_1_1_0[8|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|5] fgcell_amp_MiM_cap_1_1_0[9|5]/vinj fgcell_amp_MiM_cap_1_1_0[9|5]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|5]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|5]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|5]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|5]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|5]/vdd fgcell_amp_MiM_cap_1_1_0[9|5]/vsrc fgcell_amp_MiM_cap_1_1_0[9|5]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|6] fgcell_amp_MiM_cap_1_1_0[0|6]/vinj fgcell_amp_MiM_cap_1_1_0[0|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|6]/vdd fgcell_amp_MiM_cap_1_1_0[0|6]/vsrc fgcell_amp_MiM_cap_1_1_0[0|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|6] fgcell_amp_MiM_cap_1_1_0[1|6]/vinj fgcell_amp_MiM_cap_1_1_0[1|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|6]/vdd fgcell_amp_MiM_cap_1_1_0[1|6]/vsrc fgcell_amp_MiM_cap_1_1_0[1|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|6] fgcell_amp_MiM_cap_1_1_0[2|6]/vinj fgcell_amp_MiM_cap_1_1_0[2|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|6]/vdd fgcell_amp_MiM_cap_1_1_0[2|6]/vsrc fgcell_amp_MiM_cap_1_1_0[2|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|6] fgcell_amp_MiM_cap_1_1_0[3|6]/vinj fgcell_amp_MiM_cap_1_1_0[3|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|6]/vdd fgcell_amp_MiM_cap_1_1_0[3|6]/vsrc fgcell_amp_MiM_cap_1_1_0[3|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|6] fgcell_amp_MiM_cap_1_1_0[4|6]/vinj fgcell_amp_MiM_cap_1_1_0[4|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|6]/vdd fgcell_amp_MiM_cap_1_1_0[4|6]/vsrc fgcell_amp_MiM_cap_1_1_0[4|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|6] fgcell_amp_MiM_cap_1_1_0[5|6]/vinj fgcell_amp_MiM_cap_1_1_0[5|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|6]/vdd fgcell_amp_MiM_cap_1_1_0[5|6]/vsrc fgcell_amp_MiM_cap_1_1_0[5|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|6] fgcell_amp_MiM_cap_1_1_0[6|6]/vinj fgcell_amp_MiM_cap_1_1_0[6|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|6]/vdd fgcell_amp_MiM_cap_1_1_0[6|6]/vsrc fgcell_amp_MiM_cap_1_1_0[6|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|6] fgcell_amp_MiM_cap_1_1_0[7|6]/vinj fgcell_amp_MiM_cap_1_1_0[7|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|6]/vdd fgcell_amp_MiM_cap_1_1_0[7|6]/vsrc fgcell_amp_MiM_cap_1_1_0[7|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|6] fgcell_amp_MiM_cap_1_1_0[8|6]/vinj fgcell_amp_MiM_cap_1_1_0[8|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|6]/vdd fgcell_amp_MiM_cap_1_1_0[8|6]/vsrc fgcell_amp_MiM_cap_1_1_0[8|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|6] fgcell_amp_MiM_cap_1_1_0[9|6]/vinj fgcell_amp_MiM_cap_1_1_0[9|6]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|6]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|6]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|6]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|6]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|6]/vdd fgcell_amp_MiM_cap_1_1_0[9|6]/vsrc fgcell_amp_MiM_cap_1_1_0[9|6]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|7] fgcell_amp_MiM_cap_1_1_0[0|7]/vinj fgcell_amp_MiM_cap_1_1_0[0|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|7]/vdd fgcell_amp_MiM_cap_1_1_0[0|7]/vsrc fgcell_amp_MiM_cap_1_1_0[0|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|7] fgcell_amp_MiM_cap_1_1_0[1|7]/vinj fgcell_amp_MiM_cap_1_1_0[1|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|7]/vdd fgcell_amp_MiM_cap_1_1_0[1|7]/vsrc fgcell_amp_MiM_cap_1_1_0[1|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|7] fgcell_amp_MiM_cap_1_1_0[2|7]/vinj fgcell_amp_MiM_cap_1_1_0[2|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|7]/vdd fgcell_amp_MiM_cap_1_1_0[2|7]/vsrc fgcell_amp_MiM_cap_1_1_0[2|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|7] fgcell_amp_MiM_cap_1_1_0[3|7]/vinj fgcell_amp_MiM_cap_1_1_0[3|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|7]/vdd fgcell_amp_MiM_cap_1_1_0[3|7]/vsrc fgcell_amp_MiM_cap_1_1_0[3|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|7] fgcell_amp_MiM_cap_1_1_0[4|7]/vinj fgcell_amp_MiM_cap_1_1_0[4|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|7]/vdd fgcell_amp_MiM_cap_1_1_0[4|7]/vsrc fgcell_amp_MiM_cap_1_1_0[4|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|7] fgcell_amp_MiM_cap_1_1_0[5|7]/vinj fgcell_amp_MiM_cap_1_1_0[5|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|7]/vdd fgcell_amp_MiM_cap_1_1_0[5|7]/vsrc fgcell_amp_MiM_cap_1_1_0[5|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|7] fgcell_amp_MiM_cap_1_1_0[6|7]/vinj fgcell_amp_MiM_cap_1_1_0[6|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|7]/vdd fgcell_amp_MiM_cap_1_1_0[6|7]/vsrc fgcell_amp_MiM_cap_1_1_0[6|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|7] fgcell_amp_MiM_cap_1_1_0[7|7]/vinj fgcell_amp_MiM_cap_1_1_0[7|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|7]/vdd fgcell_amp_MiM_cap_1_1_0[7|7]/vsrc fgcell_amp_MiM_cap_1_1_0[7|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|7] fgcell_amp_MiM_cap_1_1_0[8|7]/vinj fgcell_amp_MiM_cap_1_1_0[8|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|7]/vdd fgcell_amp_MiM_cap_1_1_0[8|7]/vsrc fgcell_amp_MiM_cap_1_1_0[8|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|7] fgcell_amp_MiM_cap_1_1_0[9|7]/vinj fgcell_amp_MiM_cap_1_1_0[9|7]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|7]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|7]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|7]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|7]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|7]/vdd fgcell_amp_MiM_cap_1_1_0[9|7]/vsrc fgcell_amp_MiM_cap_1_1_0[9|7]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|8] fgcell_amp_MiM_cap_1_1_0[0|8]/vinj fgcell_amp_MiM_cap_1_1_0[0|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|8]/vdd fgcell_amp_MiM_cap_1_1_0[0|8]/vsrc fgcell_amp_MiM_cap_1_1_0[0|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|8] fgcell_amp_MiM_cap_1_1_0[1|8]/vinj fgcell_amp_MiM_cap_1_1_0[1|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|8]/vdd fgcell_amp_MiM_cap_1_1_0[1|8]/vsrc fgcell_amp_MiM_cap_1_1_0[1|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|8] fgcell_amp_MiM_cap_1_1_0[2|8]/vinj fgcell_amp_MiM_cap_1_1_0[2|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|8]/vdd fgcell_amp_MiM_cap_1_1_0[2|8]/vsrc fgcell_amp_MiM_cap_1_1_0[2|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|8] fgcell_amp_MiM_cap_1_1_0[3|8]/vinj fgcell_amp_MiM_cap_1_1_0[3|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|8]/vdd fgcell_amp_MiM_cap_1_1_0[3|8]/vsrc fgcell_amp_MiM_cap_1_1_0[3|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|8] fgcell_amp_MiM_cap_1_1_0[4|8]/vinj fgcell_amp_MiM_cap_1_1_0[4|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|8]/vdd fgcell_amp_MiM_cap_1_1_0[4|8]/vsrc fgcell_amp_MiM_cap_1_1_0[4|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|8] fgcell_amp_MiM_cap_1_1_0[5|8]/vinj fgcell_amp_MiM_cap_1_1_0[5|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|8]/vdd fgcell_amp_MiM_cap_1_1_0[5|8]/vsrc fgcell_amp_MiM_cap_1_1_0[5|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|8] fgcell_amp_MiM_cap_1_1_0[6|8]/vinj fgcell_amp_MiM_cap_1_1_0[6|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|8]/vdd fgcell_amp_MiM_cap_1_1_0[6|8]/vsrc fgcell_amp_MiM_cap_1_1_0[6|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|8] fgcell_amp_MiM_cap_1_1_0[7|8]/vinj fgcell_amp_MiM_cap_1_1_0[7|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|8]/vdd fgcell_amp_MiM_cap_1_1_0[7|8]/vsrc fgcell_amp_MiM_cap_1_1_0[7|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|8] fgcell_amp_MiM_cap_1_1_0[8|8]/vinj fgcell_amp_MiM_cap_1_1_0[8|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|8]/vdd fgcell_amp_MiM_cap_1_1_0[8|8]/vsrc fgcell_amp_MiM_cap_1_1_0[8|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|8] fgcell_amp_MiM_cap_1_1_0[9|8]/vinj fgcell_amp_MiM_cap_1_1_0[9|8]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|8]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|8]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|8]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|8]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|8]/vdd fgcell_amp_MiM_cap_1_1_0[9|8]/vsrc fgcell_amp_MiM_cap_1_1_0[9|8]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[0|9] fgcell_amp_MiM_cap_1_1_0[0|9]/vinj fgcell_amp_MiM_cap_1_1_0[0|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[0|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[0|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[0|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[0|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[0|9]/vdd fgcell_amp_MiM_cap_1_1_0[0|9]/vsrc fgcell_amp_MiM_cap_1_1_0[0|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[1|9] fgcell_amp_MiM_cap_1_1_0[1|9]/vinj fgcell_amp_MiM_cap_1_1_0[1|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[1|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[1|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[1|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[1|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[1|9]/vdd fgcell_amp_MiM_cap_1_1_0[1|9]/vsrc fgcell_amp_MiM_cap_1_1_0[1|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[2|9] fgcell_amp_MiM_cap_1_1_0[2|9]/vinj fgcell_amp_MiM_cap_1_1_0[2|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[2|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[2|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[2|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[2|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[2|9]/vdd fgcell_amp_MiM_cap_1_1_0[2|9]/vsrc fgcell_amp_MiM_cap_1_1_0[2|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[3|9] fgcell_amp_MiM_cap_1_1_0[3|9]/vinj fgcell_amp_MiM_cap_1_1_0[3|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[3|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[3|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[3|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[3|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[3|9]/vdd fgcell_amp_MiM_cap_1_1_0[3|9]/vsrc fgcell_amp_MiM_cap_1_1_0[3|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[4|9] fgcell_amp_MiM_cap_1_1_0[4|9]/vinj fgcell_amp_MiM_cap_1_1_0[4|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[4|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[4|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[4|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[4|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[4|9]/vdd fgcell_amp_MiM_cap_1_1_0[4|9]/vsrc fgcell_amp_MiM_cap_1_1_0[4|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[5|9] fgcell_amp_MiM_cap_1_1_0[5|9]/vinj fgcell_amp_MiM_cap_1_1_0[5|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[5|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[5|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[5|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[5|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[5|9]/vdd fgcell_amp_MiM_cap_1_1_0[5|9]/vsrc fgcell_amp_MiM_cap_1_1_0[5|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[6|9] fgcell_amp_MiM_cap_1_1_0[6|9]/vinj fgcell_amp_MiM_cap_1_1_0[6|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[6|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[6|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[6|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[6|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[6|9]/vdd fgcell_amp_MiM_cap_1_1_0[6|9]/vsrc fgcell_amp_MiM_cap_1_1_0[6|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[7|9] fgcell_amp_MiM_cap_1_1_0[7|9]/vinj fgcell_amp_MiM_cap_1_1_0[7|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[7|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[7|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[7|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[7|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[7|9]/vdd fgcell_amp_MiM_cap_1_1_0[7|9]/vsrc fgcell_amp_MiM_cap_1_1_0[7|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[8|9] fgcell_amp_MiM_cap_1_1_0[8|9]/vinj fgcell_amp_MiM_cap_1_1_0[8|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[8|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[8|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[8|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[8|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[8|9]/vdd fgcell_amp_MiM_cap_1_1_0[8|9]/vsrc fgcell_amp_MiM_cap_1_1_0[8|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
Xfgcell_amp_MiM_cap_1_1_0[9|9] fgcell_amp_MiM_cap_1_1_0[9|9]/vinj fgcell_amp_MiM_cap_1_1_0[9|9]/vtun
+ fgcell_amp_MiM_cap_1_1_0[9|9]/x1/tg5v0_0/vout fgcell_amp_MiM_cap_1_1_0[9|9]/row_en
+ fgcell_amp_MiM_cap_1_1_0[9|9]/x1/x1/vctrl fgcell_amp_MiM_cap_1_1_0[9|9]/x1/x2/vb
+ fgcell_amp_MiM_cap_1_1_0[9|9]/vdd fgcell_amp_MiM_cap_1_1_0[9|9]/vsrc fgcell_amp_MiM_cap_1_1_0[9|9]/row_en_b
+ VSUBS fgcell_amp_MiM_cap_1_1
.ends

.subckt array_core VPWR a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] VTUN VINJ VCTRL
+ VSRC c[8] c[11] c[14] c[2] c[7] c[5] c[10] c[13] c[6] c[4] c[1] c[9] r_vout c[12]
+ VOUT0 c[15] c[0] VGND c[3]
Xarray_column_decode_0 a[3] a[2] a[1] a[0] c[15] c[14] c[13] c[12] c[11] c[10] c[9]
+ c[7] c[6] c[5] c[4] c[3] c[2] c[1] c[0] c[8] VGND VPWR array_column_decode
Xarray_core_block5_0 tg5v0_1[3]/vin VTUN tg5v0_1[7]/vin array_core_block_routing_0/vctrl
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ tg5v0_1[4]/vin array_core_block_routing_0/VSRC tg5v0_1[8]/vin array_core_block_routing_0/vb
+ VTUN r_row_en[23] array_core_block_routing_0/vb array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vb tg5v0_1[1]/vin array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ r_row_en[20] tg5v0_1[2]/vin array_core_block_routing_0/vb r_row_en[29] array_core_block_routing_0/vb
+ r_row_en[23] VTUN array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC r_row_en[23] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ tg5v0_1[5]/vin array_core_block_routing_0/vb tg5v0_1[9]/vin array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vb VTUN array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ array_core_block_routing_0/VSRC VTUN tg5v0_1[6]/vin array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vb r_row_en[20] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ r_row_en[29] r_row_en[23] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ array_core_block_routing_0/vb tg5v0_1[7]/vin array_core_block_routing_0/vb array_core_block_routing_0/VSRC
+ tg5v0_1[3]/vin array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ array_core_block_routing_0/VSRC r_row_en[20] VTUN array_core_block_routing_0/vctrl
+ r_row_en[20] r_row_en[29] tg5v0_1[0]/vin tg5v0_1[4]/vin tg5v0_1[1]/vin tg5v0_1[5]/vin
+ VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ r_row_en[20] r_row_en[29] r_row_en[23] VTUN array_core_block_routing_0/vb array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj array_core_block_routing_0/VSRC array_core_block_routing_0/vb
+ array_core_block_routing_0/vb r_row_en[20] tg5v0_1[8]/vin r_row_en[29] array_core_block_routing_0/VSRC
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vb array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj tg5v0_1[9]/vin array_core_block_routing_0/vinj r_row_en[23]
+ VTUN VTUN array_core_block_routing_0/VSRC r_row_en[20] array_core_block_routing_0/vinj
+ r_row_en[29] tg5v0_1[2]/vin tg5v0_1[6]/vin VTUN array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj tg5v0_1[3]/vin array_core_block_routing_0/vinj
+ tg5v0_1[7]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vb array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vb r_row_en[20] r_row_en[29] array_core_block_routing_0/vinj
+ tg5v0_1[4]/vin r_row_en[26] array_core_block_routing_0/vb VTUN array_core_block_routing_0/vb
+ tg5v0_1[0]/vin array_core_block_routing_0/VSRC VTUN VTUN array_core_block_routing_0/vb
+ tg5v0_1[1]/vin array_core_block_routing_0/vb array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl
+ tg5v0_1[2]/vin r_row_en[26] array_core_block_routing_0/vinj r_row_en[20] r_row_en[29]
+ array_core_block_routing_0/VSRC array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vb array_core_block_routing_0/VSRC tg5v0_1[8]/vin array_core_block_routing_0/vb
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ tg5v0_1[5]/vin array_core_block_routing_0/vinj VTUN array_core_block_routing_0/VSRC
+ tg5v0_1[9]/vin array_core_block_routing_0/vb array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj array_core_block_routing_0/vb array_core_block_routing_0/vb
+ array_core_block_routing_0/vctrl tg5v0_1[6]/vin array_core_block_routing_0/VSRC
+ VTUN array_core_block_routing_0/vctrl array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ VTUN array_core_block_routing_0/vinj VTUN tg5v0_1[3]/vin array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl tg5v0_1[0]/vin
+ VTUN tg5v0_1[4]/vin r_row_en[22] array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/VSRC tg5v0_1[1]/vin array_core_block_routing_0/vb
+ array_core_block_routing_0/vctrl VTUN array_core_block_routing_0/vb array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vinj array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb array_core_block_routing_0/VSRC array_core_block_routing_0/vb
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj r_row_en[26] VTUN tg5v0_1[7]/vin array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj VTUN array_core_block_routing_0/vb array_core_block_routing_0/vb
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl tg5v0_1[8]/vin
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj VTUN r_row_en[22]
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj tg5v0_1[9]/vin array_core_block_routing_0/vinj VTUN
+ array_core_block_routing_0/vinj VTUN tg5v0_1[5]/vin array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vinj r_row_en[22]
+ array_core_block_routing_0/VSRC tg5v0_1[2]/vin array_core_block_routing_0/vb array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl tg5v0_1[6]/vin array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/vinj tg5v0_1[3]/vin array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj tg5v0_1[7]/vin array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb VTUN r_row_en[22] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb tg5v0_1[0]/vin array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ array_core_block_routing_0/VSRC VTUN array_core_block_routing_0/vinj tg5v0_1[1]/vin
+ array_core_block_routing_0/vinj r_row_en[28] VTUN r_row_en[22] array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj VTUN VTUN array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ r_row_en[22] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC tg5v0_1[4]/vin
+ array_core_block_routing_0/vb tg5v0_1[8]/vin array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC VTUN r_row_en_b[21] array_core_block_routing_0/vb
+ VTUN array_core_block_routing_0/vb VTUN tg5v0_1[5]/vin tg5v0_1[9]/vin array_core_block_routing_0/VSRC
+ r_row_en[28] r_row_en[22] r_row_en_b[23] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ r_row_en[26] tg5v0_1[6]/vin VTUN array_core_block_routing_0/vctrl tg5v0_1[2]/vin
+ array_core_block_routing_0/VSRC r_row_en_b[20] r_row_en_b[26] array_core_block_routing_0/vinj
+ r_row_en[28] VTUN r_row_en[22] tg5v0_1[3]/vin VTUN array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj r_row_en[26] r_row_en_b[22] r_row_en_b[28] tg5v0_1[0]/vin
+ array_core_block_routing_0/vctrl tg5v0_1[4]/vin array_core_block_routing_0/vb array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vb VTUN r_row_en_b[24] array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vb r_row_en[28] array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC r_row_en[22] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ VTUN array_core_block_routing_0/vb r_row_en[26] array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vinj array_core_block_routing_0/VSRC r_row_en_b[20] array_core_block_routing_0/vb
+ array_core_block_routing_0/vb array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ r_row_en[25] tg5v0_1[7]/vin r_row_en[29] r_row_en[28] array_core_block_routing_0/vinj
+ r_row_en_b[29] array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vinj array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ VTUN r_row_en_b[22] array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ tg5v0_1[8]/vin array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC VTUN array_core_block_routing_0/vctrl VTUN array_core_block_routing_0/vctrl
+ r_row_en_b[25] r_row_en[28] array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vb tg5v0_1[1]/vin array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vb tg5v0_1[5]/vin array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/vctrl VTUN VTUN r_row_en_b[21] r_row_en_b[27] array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vinj tg5v0_1[2]/vin array_core_block_routing_0/vinj tg5v0_1[6]/vin
+ r_row_en[24] array_core_block_routing_0/vinj array_core_block_routing_0/vb array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vb array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl r_row_en_b[23] r_row_en[28] r_row_en_b[29] array_core_block_routing_0/vctrl
+ r_row_en_b[22] VTUN array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ tg5v0_1[3]/vin r_row_en_b[28] VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj r_row_en_b[24] r_row_en_b[26] r_row_en[24] VTUN
+ array_core_block_routing_0/vinj array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ r_row_en_b[25] array_core_block_routing_0/vctrl r_row_en[25] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj VTUN tg5v0_1[0]/vin array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl tg5v0_1[9]/vin array_core_block_routing_0/vinj
+ r_row_en_b[28] array_core_block_routing_0/vinj VTUN array_core_block_routing_0/vctrl
+ r_row_en_b[27] VTUN tg5v0_1[1]/vin VTUN array_core_block_routing_0/VSRC r_row_en[24]
+ array_core_block_routing_0/vb r_row_en_b[23] array_core_block_routing_0/vb r_row_en_b[29]
+ r_row_en[25] array_core_block_routing_0/vinj array_core_block_routing_0/vb r_row_en[28]
+ array_core_block_routing_0/vctrl r_row_en_b[25] array_core_block_routing_0/vctrl
+ VTUN r_row_en[22] array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ tg5v0_1[7]/vin array_core_block_routing_0/vb array_core_block_routing_0/VSRC array_core_block_routing_0/vb
+ r_row_en_b[20] array_core_block_routing_0/vb r_row_en_b[26] r_row_en[24] VTUN array_core_block_routing_0/vinj
+ tg5v0_1[4]/vin tg5v0_1[8]/vin VTUN array_core_block_routing_0/VSRC r_row_en_b[22]
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj r_row_en_b[21] array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vctrl tg5v0_1[5]/vin
+ array_core_block_routing_0/vinj tg5v0_1[9]/vin VTUN r_row_en_b[24] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj r_row_en[24] r_row_en_b[23] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj r_row_en_b[25] array_core_block_routing_0/vinj VTUN
+ tg5v0_1[2]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ r_row_en_b[21] array_core_block_routing_0/VSRC VTUN r_row_en_b[27] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj r_row_en_b[20] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ r_row_en_b[26] array_core_block_routing_0/vinj array_core_block_routing_0/vb tg5v0_1[3]/vin
+ r_row_en[21] array_core_block_routing_0/vb r_row_en[24] r_row_en_b[23] VTUN r_row_en[25]
+ r_row_en_b[29] array_core_block_routing_0/vinj array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ r_row_en_b[22] tg5v0_1[0]/vin r_row_en_b[28] array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/vinj r_row_en_b[24] VTUN r_row_en[24] array_core_block_routing_0/vb
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vinj r_row_en[25] tg5v0_1[6]/vin
+ VTUN r_row_en[25] array_core_block_routing_0/VSRC r_row_en_b[27] r_row_en_b[21]
+ array_core_block_routing_0/vinj array_core_block_routing_0/VSRC r_row_en_b[20] array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC tg5v0_1[7]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb r_row_en[21] array_core_block_routing_0/vinj r_row_en[26]
+ r_row_en_b[29] array_core_block_routing_0/vinj r_row_en[24] r_row_en_b[23] VTUN
+ array_core_block_routing_0/VSRC tg5v0_1[8]/vin array_core_block_routing_0/vinj VTUN
+ r_row_en[25] array_core_block_routing_0/vb array_core_block_routing_0/vb tg5v0_1[4]/vin
+ r_row_en[29] r_row_en_b[20] array_core_block_routing_0/vinj VTUN array_core_block_routing_0/VSRC
+ r_row_en_b[26] array_core_block_routing_0/vinj r_row_en[21] r_row_en_b[25] tg5v0_1[1]/vin
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl r_row_en[26] array_core_block_routing_0/vb
+ tg5v0_1[5]/vin array_core_block_routing_0/vb VTUN array_core_block_routing_0/vinj
+ r_row_en_b[22] array_core_block_routing_0/vinj VTUN r_row_en_b[28] VTUN r_row_en_b[21]
+ r_row_en_b[27] tg5v0_1[2]/vin r_row_en[25] tg5v0_1[6]/vin array_core_block_routing_0/VSRC
+ r_row_en_b[24] array_core_block_routing_0/vinj VTUN array_core_block_routing_0/VSRC
+ array_core_block_routing_0/VSRC r_row_en[21] r_row_en_b[23] r_row_en_b[29] array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj r_row_en_b[25]
+ array_core_block_routing_0/vinj r_row_en[24] array_core_block_routing_0/vinj r_row_en[28]
+ VTUN array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vinj r_row_en_b[27] r_row_en_b[26]
+ tg5v0_1[0]/vin array_core_block_routing_0/vinj r_row_en[27] array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj r_row_en[21] tg5v0_1[9]/vin array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl r_row_en_b[29]
+ array_core_block_routing_0/vb array_core_block_routing_0/vb r_row_en_b[28] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/vb
+ array_core_block_routing_0/vb VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj r_row_en_b[24]
+ array_core_block_routing_0/vb array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ r_row_en[27] array_core_block_routing_0/VSRC array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ VTUN r_row_en[21] array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ r_row_en_b[25] array_core_block_routing_0/vctrl array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj tg5v0_1[3]/vin VTUN array_core_block_routing_0/vinj
+ tg5v0_1[7]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ array_core_block_routing_0/vctrl VTUN array_core_block_routing_0/vinj VTUN array_core_block_routing_0/VSRC
+ r_row_en_b[21] r_row_en_b[27] array_core_block_routing_0/vinj array_core_block_routing_0/vctrl
+ r_row_en_b[20] array_core_block_routing_0/vinj tg5v0_1[4]/vin tg5v0_1[8]/vin r_row_en[27]
+ VTUN array_core_block_routing_0/VSRC r_row_en[21] r_row_en_b[23] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj r_row_en_b[22] tg5v0_1[5]/vin array_core_block_routing_0/vinj
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vctrl VTUN tg5v0_1[1]/vin
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj r_row_en_b[24]
+ array_core_block_routing_0/vinj r_row_en_b[26] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ r_row_en_b[25] r_row_en[27] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ VTUN array_core_block_routing_0/VSRC tg5v0_1[2]/vin r_row_en[21] array_core_block_routing_0/vb
+ VTUN r_row_en_b[22] r_row_en_b[28] array_core_block_routing_0/vctrl r_row_en_b[21]
+ array_core_block_routing_0/vctrl array_core_block_routing_0/vinj r_row_en_b[27]
+ array_core_block_routing_0/vinj tg5v0_1[3]/vin r_row_en[21] array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vb array_core_block_routing_0/vb array_core_block_routing_0/vctrl
+ r_row_en_b[24] r_row_en_b[23] VTUN r_row_en[27] r_row_en_b[29] array_core_block_routing_0/vinj
+ r_row_en[21] VTUN array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj VTUN tg5v0_1[9]/vin array_core_block_routing_0/VSRC
+ VTUN array_core_block_routing_0/vctrl VTUN array_core_block_routing_0/vinj VTUN
+ r_row_en_b[20] tg5v0_1[6]/vin r_row_en[27] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj r_row_en[20] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vb VTUN array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ r_row_en_b[28] r_row_en_b[22] array_core_block_routing_0/vinj VTUN r_row_en_b[21]
+ array_core_block_routing_0/vinj tg5v0_1[7]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vb array_core_block_routing_0/vinj
+ array_core_block_routing_0/vb r_row_en_b[24] array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ r_row_en_b[25] r_row_en[27] array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj VTUN tg5v0_1[0]/vin array_core_block_routing_0/vb
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj tg5v0_1[4]/vin array_core_block_routing_0/vb
+ array_core_block_routing_0/VSRC array_core_block_routing_0/vinj array_core_block_routing_0/vinj
+ r_row_en[24] array_core_block_routing_0/vinj r_row_en_b[21] r_row_en_b[27] r_row_en_b[20]
+ array_core_block_routing_0/vinj VTUN tg5v0_1[1]/vin r_row_en_b[26] array_core_block_routing_0/vinj
+ tg5v0_1[5]/vin r_row_en[23] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj r_row_en_b[23] r_row_en_b[29]
+ r_row_en[27] array_core_block_routing_0/VSRC r_row_en_b[22] array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/VSRC r_row_en_b[28] tg5v0_1[2]/vin array_core_block_routing_0/vinj
+ VTUN array_core_block_routing_0/vinj array_core_block_routing_0/vinj VTUN array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj r_row_en_b[24] array_core_block_routing_0/vinj array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj r_row_en_b[26] r_row_en[23] array_core_block_routing_0/vinj
+ array_core_block_routing_0/vinj VTUN array_core_block_routing_0/vinj r_row_en_b[25]
+ VTUN r_row_en[25] r_row_en[27] array_core_block_routing_0/VSRC array_core_block_routing_0/vinj
+ tg5v0_1[8]/vin array_core_block_routing_0/VSRC array_core_block_routing_0/vb VTUN
+ r_row_en_b[28] array_core_block_routing_0/vinj array_core_block_routing_0/vb r_row_en_b[27]
+ array_core_block_routing_0/vb tg5v0_1[0]/vin array_core_block_routing_0/vinj array_core_block_routing_0/vb
+ r_row_en[26] tg5v0_1[9]/vin array_core_block_routing_0/VSRC r_row_en[28] VTUN array_core_block_routing_0/VSRC
+ array_core_block_routing_0/vinj array_core_block_routing_0/vinj r_row_en[23] array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC r_row_en_b[29] array_core_block_routing_0/vb r_row_en[27]
+ array_core_block_routing_0/vctrl r_row_en[25] array_core_block_routing_0/vb VTUN
+ array_core_block_routing_0/vinj VGND VTUN array_core_block_routing_0/VSRC tg5v0_1[6]/vin
+ r_row_en_b[20] r_row_en[26] array_core_block_routing_0/VSRC r_row_en_b[26] array_core_block_routing_0/vinj
+ array_core_block_routing_0/VSRC r_row_en[23] array_core_block5
Xarray_row_decode_0 a[8] a[7] a[6] a[5] a[4] r_w[31] r_w[30] r_w[29] r_w[28] r_w[27]
+ r_w[26] r_w[25] r_w[24] r_w[23] r_w[22] r_w[21] r_w[20] r_w[19] r_w[18] r_w[17]
+ r_w[16] r_w[15] r_w[14] r_w[13] r_w[12] r_w[11] r_w[10] r_w[9] r_w[8] r_w[7] r_w[6]
+ r_w[5] r_w[4] r_w[3] r_w[2] r_w[1] r_w[0] VGND VPWR array_row_decode
Xarray_row_decode_1 a[8] a[7] a[6] a[5] a[4] l_w[31] l_w[30] l_w[29] l_w[28] l_w[27]
+ l_w[26] l_w[25] l_w[24] l_w[23] l_w[22] l_w[21] l_w[20] l_w[19] l_w[18] l_w[17]
+ l_w[16] l_w[15] l_w[14] l_w[13] l_w[12] l_w[11] l_w[10] l_w[9] l_w[8] l_w[7] l_w[6]
+ l_w[5] l_w[4] l_w[3] l_w[2] l_w[1] l_w[0] VGND VPWR array_row_decode
Xarray_core_block1_0 VTUN VSRC VSRC l_row_en[10] l_row_en[14] tg5v0_0[6]/vin vb l_row_en[13]
+ VCTRL VCTRL VCTRL l_row_en[16] vb VINJ tg5v0_0[0]/vin VTUN l_row_en[19] l_row_en[15]
+ VTUN VSRC tg5v0_0[0]/vin VCTRL VCTRL VCTRL tg5v0_0[5]/vin vb VINJ tg5v0_0[5]/vin
+ vb VSRC VSRC VSRC VINJ vb tg5v0_0[4]/vin vb VTUN VINJ VSRC VSRC l_row_en[10] VSRC
+ VSRC VINJ l_row_en[13] tg5v0_0[9]/vin VCTRL VCTRL l_row_en[12] vb l_row_en[15] VINJ
+ tg5v0_0[3]/vin vb VTUN VSRC VINJ VSRC l_row_en[17] tg5v0_0[3]/vin VCTRL VCTRL VCTRL
+ VCTRL VSRC tg5v0_0[8]/vin vb tg5v0_0[8]/vin VINJ vb VTUN VCTRL VCTRL VSRC VSRC tg5v0_0[2]/vin
+ vb tg5v0_0[7]/vin vb l_row_en[10] VSRC VSRC tg5v0_0[1]/vin l_row_en[12] VINJ tg5v0_0[1]/vin
+ l_row_en[15] vb l_row_en[14] tg5v0_0[6]/vin vb VTUN VSRC VCTRL VCTRL l_row_en[17]
+ VCTRL VSRC tg5v0_0[6]/vin l_row_en[19] VINJ VINJ tg5v0_0[0]/vin VINJ vb VCTRL VCTRL
+ VCTRL VSRC vb VTUN tg5v0_0[5]/vin VINJ VINJ VINJ vb VSRC VSRC l_row_en[12] tg5v0_0[4]/vin
+ vb VINJ l_row_en[14] VTUN VINJ l_row_en[17] l_row_en[13] VCTRL VCTRL VCTRL tg5v0_0[9]/vin
+ VSRC l_row_en[16] VSRC l_row_en[19] tg5v0_0[3]/vin vb VINJ VINJ tg5v0_0[3]/vin VCTRL
+ VCTRL VCTRL VINJ VTUN VINJ vb tg5v0_0[8]/vin VTUN VSRC VSRC tg5v0_0[8]/vin VINJ
+ vb VINJ VINJ VINJ tg5v0_0[2]/vin VTUN VTUN VSRC vb VSRC tg5v0_0[7]/vin l_row_en[10]
+ vb VINJ l_row_en[13] VCTRL VCTRL VCTRL VTUN VINJ tg5v0_0[1]/vin VTUN l_row_en[16]
+ vb VSRC tg5v0_0[1]/vin l_row_en[15] tg5v0_0[6]/vin VINJ VCTRL VCTRL VCTRL VCTRL
+ VINJ l_row_en[11] tg5v0_0[6]/vin vb VINJ VINJ VINJ VTUN VTUN VSRC VSRC vb VSRC tg5v0_0[0]/vin
+ VCTRL VINJ VINJ vb VINJ tg5v0_0[5]/vin VTUN VINJ VINJ VTUN VSRC vb VSRC VSRC l_row_en[10]
+ VINJ l_row_en[13] VCTRL l_row_en[12] tg5v0_0[4]/vin vb VINJ VINJ VINJ VTUN l_row_en[15]
+ VSRC VSRC vb tg5v0_0[4]/vin VSRC l_row_en[17] tg5v0_0[9]/vin VCTRL VCTRL VCTRL VTUN
+ tg5v0_0[9]/vin vb VINJ VINJ VTUN VTUN VSRC VINJ VINJ vb VSRC VINJ tg5v0_0[3]/vin
+ VCTRL VCTRL l_row_en[18] VINJ VTUN VTUN VINJ tg5v0_0[8]/vin vb VINJ VTUN VTUN VSRC
+ VSRC vb tg5v0_0[2]/vin l_row_en[10] VINJ l_row_en[12] VTUN VINJ VINJ tg5v0_0[7]/vin
+ l_row_en[15] vb VSRC l_row_en[18] VTUN l_row_en[14] VSRC VINJ vb VSRC l_row_en[17]
+ VCTRL VCTRL tg5v0_0[1]/vin VCTRL l_row_en[16] VINJ tg5v0_0[1]/vin l_row_en[19] VINJ
+ VTUN tg5v0_0[6]/vin VTUN VSRC VCTRL VCTRL VCTRL VINJ l_row_en_b[18] VSRC VSRC vb
+ VINJ tg5v0_0[6]/vin VTUN l_row_en_b[11] VINJ VINJ tg5v0_0[0]/vin l_row_en_b[18]
+ vb VINJ VTUN VINJ VSRC VTUN VSRC VSRC tg5v0_0[5]/vin VTUN l_row_en_b[15] vb VINJ
+ l_row_en[14] VTUN VTUN VSRC VINJ VINJ l_row_en[13] VCTRL VCTRL VCTRL VCTRL vb VSRC
+ VINJ l_row_en[16] l_row_en_b[15] tg5v0_0[4]/vin l_row_en[19] tg5v0_0[4]/vin VTUN
+ VTUN l_row_en_b[12] vb VINJ VCTRL VCTRL VCTRL VCTRL VTUN tg5v0_0[9]/vin VSRC VINJ
+ vb l_row_en_b[19] VSRC tg5v0_0[9]/vin vb l_row_en_b[12] VTUN VINJ VINJ tg5v0_0[3]/vin
+ l_row_en_b[19] vb VSRC VTUN VINJ VSRC vb VINJ l_row_en_b[16] tg5v0_0[8]/vin vb VINJ
+ VINJ tg5v0_0[2]/vin l_row_en[10] l_row_en_b[16] VTUN l_row_en[11] vb VSRC l_row_en[13]
+ VCTRL VCTRL VTUN VINJ VSRC tg5v0_0[2]/vin l_row_en[16] vb VTUN VINJ VINJ l_row_en_b[13]
+ VINJ tg5v0_0[7]/vin l_row_en[15] vb VSRC VINJ VINJ l_row_en_b[17] tg5v0_0[7]/vin
+ VCTRL VCTRL VCTRL l_row_en_b[13] VTUN vb VSRC VTUN tg5v0_0[1]/vin l_row_en_b[14]
+ l_row_en[11] VSRC vb l_row_en_b[10] VINJ vb VCTRL VINJ VINJ VINJ l_row_en_b[17]
+ VTUN l_row_en_b[14] tg5v0_0[6]/vin VTUN VTUN l_row_en_b[10] vb VSRC VINJ VSRC VINJ
+ tg5v0_0[0]/vin vb VINJ VINJ l_row_en_b[17] VINJ vb l_row_en[10] VINJ VINJ VINJ l_row_en[13]
+ VCTRL l_row_en_b[11] VTUN tg5v0_0[5]/vin l_row_en[12] vb VSRC l_row_en_b[18] l_row_en[15]
+ VSRC l_row_en_b[14] vb l_row_en_b[11] l_row_en[14] vb VTUN VCTRL VINJ VINJ l_row_en[17]
+ VCTRL VCTRL VINJ VINJ VTUN VTUN l_row_en[18] VINJ l_row_en_b[14] tg5v0_0[4]/vin
+ VTUN l_row_en[19] vb VSRC VINJ l_row_en_b[15] tg5v0_0[4]/vin vb l_row_en_b[11] VINJ
+ VCTRL VCTRL tg5v0_0[9]/vin vb VINJ VINJ l_row_en_b[18] VTUN VINJ l_row_en_b[15]
+ tg5v0_0[9]/vin VTUN l_row_en_b[11] VTUN VINJ l_row_en[18] vb VTUN l_row_en_b[12]
+ VINJ tg5v0_0[3]/vin vb VINJ l_row_en_b[19] vb VINJ VINJ l_row_en_b[15] VINJ VINJ
+ l_row_en_b[12] l_row_en[12] VTUN VTUN tg5v0_0[8]/vin VSRC VINJ l_row_en[11] VSRC
+ l_row_en_b[19] l_row_en[14] l_row_en_b[15] tg5v0_0[2]/vin vb VINJ l_row_en[17] l_row_en[18]
+ VCTRL VCTRL VCTRL VCTRL VINJ tg5v0_0[2]/vin l_row_en_b[16] vb VINJ l_row_en_b[18]
+ l_row_en[16] VTUN VINJ l_row_en_b[12] VTUN VINJ l_row_en[19] VTUN tg5v0_0[7]/vin
+ vb VSRC VINJ l_row_en_b[19] VSRC VINJ VINJ tg5v0_0[7]/vin l_row_en_b[16] VCTRL VCTRL
+ VCTRL VCTRL VINJ l_row_en_b[12] VINJ l_row_en_b[13] vb VTUN VINJ tg5v0_0[1]/vin
+ l_row_en_b[19] VINJ VINJ VTUN VTUN vb VSRC l_row_en_b[16] VSRC l_row_en_b[13] vb
+ VINJ tg5v0_0[6]/vin VTUN VINJ VTUN VTUN tg5v0_0[0]/vin l_row_en_b[16] VINJ VINJ
+ VINJ l_row_en[11] VTUN VTUN VSRC tg5v0_0[0]/vin vb l_row_en[14] l_row_en_b[10] l_row_en[13]
+ VCTRL VCTRL VCTRL vb tg5v0_0[5]/vin l_row_en[16] vb VINJ VINJ l_row_en_b[17] tg5v0_0[5]/vin
+ VINJ l_row_en[19] VTUN VINJ VINJ l_row_en_b[13] VINJ l_row_en[18] l_row_en_b[10]
+ VTUN VTUN vb VSRC VCTRL VCTRL VCTRL l_row_en_b[17] vb VINJ VINJ l_row_en_b[13] vb
+ l_row_en_b[14] VINJ tg5v0_0[4]/vin VTUN VINJ VINJ l_row_en_b[10] VTUN VSRC VINJ
+ l_row_en[11] VTUN VSRC vb VSRC l_row_en_b[17] l_row_en_b[14] vb tg5v0_0[9]/vin l_row_en_b[10]
+ vb VINJ l_row_en[11] l_row_en_b[11] VINJ VINJ l_row_en_b[17] tg5v0_0[3]/vin VTUN
+ VSRC l_row_en[10] VTUN l_row_en_b[18] vb VSRC VINJ l_row_en[13] VCTRL VCTRL VSRC
+ l_row_en_b[14] l_row_en[11] tg5v0_0[8]/vin l_row_en[16] l_row_en[12] l_row_en_b[11]
+ vb l_row_en[15] VINJ vb l_row_en_b[18] VINJ l_row_en[18] tg5v0_0[2]/vin VTUN l_row_en_b[14]
+ VINJ l_row_en[17] VCTRL VCTRL VCTRL VTUN VSRC l_row_en_b[15] VSRC tg5v0_0[2]/vin
+ vb VINJ l_row_en_b[11] vb VINJ tg5v0_0[7]/vin l_row_en_b[18] l_row_en[11] vb l_row_en_b[15]
+ VTUN VINJ VINJ tg5v0_0[7]/vin VCTRL VINJ l_row_en_b[11] VTUN VINJ VSRC VINJ l_row_en_b[12]
+ vb VTUN VSRC VINJ tg5v0_0[1]/vin l_row_en_b[18] vb l_row_en_b[19] VINJ l_row_en_b[15]
+ vb VTUN VINJ l_row_en[10] l_row_en_b[12] VINJ tg5v0_0[6]/vin VTUN VINJ l_row_en[18]
+ VCTRL VSRC l_row_en_b[19] VSRC tg5v0_0[0]/vin l_row_en[12] vb VTUN l_row_en_b[15]
+ VINJ l_row_en[15] vb VINJ VINJ tg5v0_0[0]/vin l_row_en[14] VINJ vb VINJ VINJ VCTRL
+ VCTRL VINJ l_row_en[17] tg5v0_0[5]/vin VCTRL VCTRL VSRC VINJ VINJ VTUN VSRC VINJ
+ l_row_en_b[16] l_row_en[19] tg5v0_0[5]/vin vb VINJ l_row_en_b[12] l_row_en[18] VINJ
+ vb VCTRL l_row_en_b[19] VCTRL VCTRL VINJ l_row_en_b[16] vb VTUN VINJ VINJ VINJ l_row_en_b[12]
+ VTUN VSRC VINJ VSRC VINJ l_row_en_b[13] l_row_en_b[19] tg5v0_0[4]/vin VINJ vb l_row_en[18]
+ VINJ l_row_en_b[16] vb VINJ VINJ l_row_en_b[13] tg5v0_0[9]/vin VTUN VINJ VSRC VSRC
+ VINJ l_row_en[12] VTUN VSRC VINJ l_row_en[11] l_row_en_b[10] tg5v0_0[3]/vin VINJ
+ l_row_en_b[16] l_row_en_b[18] l_row_en[14] l_row_en_b[17] VINJ l_row_en[17] tg5v0_0[3]/vin
+ VCTRL VCTRL VCTRL l_row_en_b[13] VINJ vb VTUN l_row_en_b[10] tg5v0_0[8]/vin l_row_en[16]
+ VSRC VINJ VINJ VSRC VINJ l_row_en[19] VTUN VSRC VINJ l_row_en_b[17] VINJ tg5v0_0[8]/vin
+ l_row_en_b[13] vb VTUN VCTRL VCTRL VCTRL l_row_en_b[14] VINJ tg5v0_0[2]/vin l_row_en_b[10]
+ VINJ VTUN VINJ VSRC VSRC VINJ l_row_en_b[17] VTUN VSRC VINJ l_row_en_b[14] tg5v0_0[7]/vin
+ VINJ VGND l_row_en_b[10] vb VTUN VINJ VINJ VINJ tg5v0_0[1]/vin l_row_en_b[11] vb
+ VTUN array_core_block1
Xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_0 VGND vb VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield m=1
Xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_1 VGND vb VGND sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield m=1
Xlsi1v8o5v0_0[0] l_w[31] l_row_en_b[31] l_row_en[31] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[1] l_w[30] l_row_en_b[30] l_row_en[30] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[2] l_w[29] l_row_en_b[29] l_row_en[29] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[3] l_w[28] l_row_en_b[28] l_row_en[28] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[4] l_w[27] l_row_en_b[27] l_row_en[27] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[5] l_w[26] l_row_en_b[26] l_row_en[26] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[6] l_w[25] l_row_en_b[25] l_row_en[25] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[7] l_w[24] l_row_en_b[24] l_row_en[24] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[8] l_w[23] l_row_en_b[23] l_row_en[23] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[9] l_w[22] l_row_en_b[22] l_row_en[22] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[10] l_w[21] l_row_en_b[21] l_row_en[21] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[11] l_w[20] l_row_en_b[20] l_row_en[20] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[12] l_w[19] l_row_en_b[19] l_row_en[19] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[13] l_w[18] l_row_en_b[18] l_row_en[18] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[14] l_w[17] l_row_en_b[17] l_row_en[17] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[15] l_w[16] l_row_en_b[16] l_row_en[16] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[16] l_w[15] l_row_en_b[15] l_row_en[15] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[17] l_w[14] l_row_en_b[14] l_row_en[14] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[18] l_w[13] l_row_en_b[13] l_row_en[13] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[19] l_w[12] l_row_en_b[12] l_row_en[12] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[20] l_w[11] l_row_en_b[11] l_row_en[11] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[21] l_w[10] l_row_en_b[10] l_row_en[10] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[22] l_w[9] l_row_en_b[9] l_row_en[9] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[23] l_w[8] l_row_en_b[8] l_row_en[8] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[24] l_w[7] l_row_en_b[7] l_row_en[7] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[25] l_w[6] l_row_en_b[6] l_row_en[6] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[26] l_w[5] l_row_en_b[5] l_row_en[5] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[27] l_w[4] l_row_en_b[4] l_row_en[4] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[28] l_w[3] l_row_en_b[3] l_row_en[3] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[29] l_w[2] l_row_en_b[2] l_row_en[2] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[30] l_w[1] l_row_en_b[1] l_row_en[1] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_0[31] l_w[0] l_row_en_b[0] l_row_en[0] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[0] r_w[31] r_row_en_b[31] r_row_en[31] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[1] r_w[30] r_row_en_b[30] r_row_en[30] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[2] r_w[29] r_row_en_b[29] r_row_en[29] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[3] r_w[28] r_row_en_b[28] r_row_en[28] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[4] r_w[27] r_row_en_b[27] r_row_en[27] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[5] r_w[26] r_row_en_b[26] r_row_en[26] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[6] r_w[25] r_row_en_b[25] r_row_en[25] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[7] r_w[24] r_row_en_b[24] r_row_en[24] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[8] r_w[23] r_row_en_b[23] r_row_en[23] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[9] r_w[22] r_row_en_b[22] r_row_en[22] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[10] r_w[21] r_row_en_b[21] r_row_en[21] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[11] r_w[20] r_row_en_b[20] r_row_en[20] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[12] r_w[19] r_row_en_b[19] r_row_en[19] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[13] r_w[18] r_row_en_b[18] r_row_en[18] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[14] r_w[17] r_row_en_b[17] r_row_en[17] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[15] r_w[16] r_row_en_b[16] r_row_en[16] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[16] r_w[15] r_row_en_b[15] r_row_en[15] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[17] r_w[14] r_row_en_b[14] r_row_en[14] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[18] r_w[13] r_row_en_b[13] r_row_en[13] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[19] r_w[12] r_row_en_b[12] r_row_en[12] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[20] r_w[11] r_row_en_b[11] r_row_en[11] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[21] r_w[10] r_row_en_b[10] r_row_en[10] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[22] r_w[9] r_row_en_b[9] r_row_en[9] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[23] r_w[8] r_row_en_b[8] r_row_en[8] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[24] r_w[7] r_row_en_b[7] r_row_en[7] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[25] r_w[6] r_row_en_b[6] r_row_en[6] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[26] r_w[5] r_row_en_b[5] r_row_en[5] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[27] r_w[4] r_row_en_b[4] r_row_en[4] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[28] r_w[3] r_row_en_b[3] r_row_en[3] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[29] r_w[2] r_row_en_b[2] r_row_en[2] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[30] r_w[1] r_row_en_b[1] r_row_en[1] VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_1[31] r_w[0] r_row_en_b[0] r_row_en[0] VPWR VINJ VGND lsi1v8o5v0
Xtg5v0_0[0] tg5v0_0[0]/vin VOUT0 tg5v0_1[0]/en tg5v0_1[0]/en_b VINJ VGND tg5v0
Xtg5v0_0[1] tg5v0_0[1]/vin VOUT0 tg5v0_1[1]/en tg5v0_1[1]/en_b VINJ VGND tg5v0
Xtg5v0_0[2] tg5v0_0[2]/vin VOUT0 tg5v0_1[2]/en tg5v0_1[2]/en_b VINJ VGND tg5v0
Xtg5v0_0[3] tg5v0_0[3]/vin VOUT0 tg5v0_1[3]/en tg5v0_1[3]/en_b VINJ VGND tg5v0
Xtg5v0_0[4] tg5v0_0[4]/vin VOUT0 tg5v0_1[4]/en tg5v0_1[4]/en_b VINJ VGND tg5v0
Xtg5v0_0[5] tg5v0_0[5]/vin VOUT0 tg5v0_1[5]/en tg5v0_1[5]/en_b VINJ VGND tg5v0
Xtg5v0_0[6] tg5v0_0[6]/vin VOUT0 tg5v0_1[6]/en tg5v0_1[6]/en_b VINJ VGND tg5v0
Xtg5v0_0[7] tg5v0_0[7]/vin VOUT0 tg5v0_1[7]/en tg5v0_1[7]/en_b VINJ VGND tg5v0
Xtg5v0_0[8] tg5v0_0[8]/vin VOUT0 tg5v0_1[8]/en tg5v0_1[8]/en_b VINJ VGND tg5v0
Xtg5v0_0[9] tg5v0_0[9]/vin VOUT0 tg5v0_1[9]/en tg5v0_1[9]/en_b VINJ VGND tg5v0
Xlsi1v8o5v0_2[0] c[15] lsi1v8o5v0_2[0]/out_b lsi1v8o5v0_2[0]/out VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[1] c[14] lsi1v8o5v0_2[1]/out_b lsi1v8o5v0_2[1]/out VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[2] c[13] lsi1v8o5v0_2[2]/out_b lsi1v8o5v0_2[2]/out VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[3] c[12] tg5v0_2/en_b tg5v0_2/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[4] c[11] tg5v0_4/en_b tg5v0_4/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[5] c[10] tg5v0_3/en_b tg5v0_3/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[6] c[9] tg5v0_1[9]/en_b tg5v0_1[9]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[7] c[8] tg5v0_1[8]/en_b tg5v0_1[8]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[8] c[7] tg5v0_1[7]/en_b tg5v0_1[7]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[9] c[6] tg5v0_1[6]/en_b tg5v0_1[6]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[10] c[5] tg5v0_1[5]/en_b tg5v0_1[5]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[11] c[4] tg5v0_1[4]/en_b tg5v0_1[4]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[12] c[3] tg5v0_1[3]/en_b tg5v0_1[3]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[13] c[2] tg5v0_1[2]/en_b tg5v0_1[2]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[14] c[1] tg5v0_1[1]/en_b tg5v0_1[1]/en VPWR VINJ VGND lsi1v8o5v0
Xlsi1v8o5v0_2[15] c[0] tg5v0_1[0]/en_b tg5v0_1[0]/en VPWR VINJ VGND lsi1v8o5v0
Xtg5v0_1[0] tg5v0_1[0]/vin r_vout tg5v0_1[0]/en tg5v0_1[0]/en_b VINJ VGND tg5v0
Xtg5v0_1[1] tg5v0_1[1]/vin r_vout tg5v0_1[1]/en tg5v0_1[1]/en_b VINJ VGND tg5v0
Xtg5v0_1[2] tg5v0_1[2]/vin r_vout tg5v0_1[2]/en tg5v0_1[2]/en_b VINJ VGND tg5v0
Xtg5v0_1[3] tg5v0_1[3]/vin r_vout tg5v0_1[3]/en tg5v0_1[3]/en_b VINJ VGND tg5v0
Xtg5v0_1[4] tg5v0_1[4]/vin r_vout tg5v0_1[4]/en tg5v0_1[4]/en_b VINJ VGND tg5v0
Xtg5v0_1[5] tg5v0_1[5]/vin r_vout tg5v0_1[5]/en tg5v0_1[5]/en_b VINJ VGND tg5v0
Xtg5v0_1[6] tg5v0_1[6]/vin r_vout tg5v0_1[6]/en tg5v0_1[6]/en_b VINJ VGND tg5v0
Xtg5v0_1[7] tg5v0_1[7]/vin r_vout tg5v0_1[7]/en tg5v0_1[7]/en_b VINJ VGND tg5v0
Xtg5v0_1[8] tg5v0_1[8]/vin r_vout tg5v0_1[8]/en tg5v0_1[8]/en_b VINJ VGND tg5v0
Xtg5v0_1[9] tg5v0_1[9]/vin r_vout tg5v0_1[9]/en tg5v0_1[9]/en_b VINJ VGND tg5v0
Xtg5v0_2 VGND VOUT0 tg5v0_2/en tg5v0_2/en_b VINJ VGND tg5v0
Xtg5v0_3 vb VOUT0 tg5v0_3/en tg5v0_3/en_b VINJ VGND tg5v0
Xtg5v0_4 VINJ VOUT0 tg5v0_4/en tg5v0_4/en_b VINJ VGND tg5v0
Xarray_core_block2_0 l_row_en[20] VTUN VSRC l_row_en[23] tg5v0_0[7]/vin VSRC VSRC
+ VCTRL VCTRL l_row_en[26] vb tg5v0_0[1]/vin vb l_row_en[28] VTUN tg5v0_0[1]/vin vb
+ VTUN VSRC VCTRL VCTRL tg5v0_0[6]/vin VCTRL VSRC vb tg5v0_0[6]/vin vb VINJ VINJ VTUN
+ vb tg5v0_0[0]/vin VCTRL VTUN VSRC VINJ VSRC vb tg5v0_0[5]/vin vb VINJ l_row_en[20]
+ vb l_row_en[23] VTUN VSRC VSRC l_row_en[22] VCTRL VINJ l_row_en[28] l_row_en[24]
+ tg5v0_0[4]/vin vb VINJ l_row_en[27] VINJ VTUN tg5v0_0[4]/vin VCTRL VCTRL VCTRL vb
+ VSRC VTUN l_row_en[29] tg5v0_0[9]/vin tg5v0_0[9]/vin VCTRL VCTRL VINJ VTUN vb VSRC
+ tg5v0_0[3]/vin VSRC vb tg5v0_0[8]/vin VTUN VINJ VINJ VTUN l_row_en[22] VSRC tg5v0_0[2]/vin
+ l_row_en[21] VSRC tg5v0_0[2]/vin l_row_en[24] VINJ tg5v0_0[7]/vin l_row_en[27] vb
+ VINJ VTUN l_row_en[26] VCTRL VCTRL VCTRL VCTRL vb VTUN tg5v0_0[7]/vin l_row_en[29]
+ VSRC VSRC tg5v0_0[1]/vin VCTRL VCTRL VCTRL VCTRL vb VINJ vb VTUN tg5v0_0[6]/vin
+ VSRC tg5v0_0[0]/vin VINJ vb VTUN vb VTUN VINJ l_row_en[21] tg5v0_0[5]/vin l_row_en[24]
+ l_row_en[23] VINJ l_row_en[26] VCTRL VCTRL VCTRL vb l_row_en[29] VTUN vb VSRC l_row_en[28]
+ tg5v0_0[4]/vin VSRC VCTRL tg5v0_0[4]/vin VCTRL VCTRL VINJ tg5v0_0[9]/vin vb VTUN
+ vb VSRC tg5v0_0[9]/vin VSRC VINJ VINJ tg5v0_0[3]/vin VINJ VINJ vb VINJ l_row_en[21]
+ vb VSRC tg5v0_0[8]/vin l_row_en[20] VSRC l_row_en[23] l_row_en[26] VCTRL VCTRL tg5v0_0[2]/vin
+ l_row_en[22] VINJ VTUN VINJ vb tg5v0_0[2]/vin l_row_en[28] VTUN VINJ vb VSRC VINJ
+ tg5v0_0[7]/vin l_row_en[27] VCTRL VCTRL VCTRL tg5v0_0[7]/vin VINJ VINJ VTUN VINJ
+ vb tg5v0_0[1]/vin VTUN VSRC VCTRL vb tg5v0_0[6]/vin VTUN VINJ VINJ VINJ vb VTUN
+ VSRC tg5v0_0[0]/vin l_row_en[20] vb VSRC VINJ VINJ tg5v0_0[0]/vin l_row_en[22] VCTRL
+ tg5v0_0[5]/vin VINJ l_row_en[24] VTUN tg5v0_0[5]/vin l_row_en[27] VSRC VINJ VCTRL
+ VCTRL VCTRL VCTRL vb VTUN VINJ l_row_en[29] l_row_en[25] vb VINJ VTUN VINJ tg5v0_0[4]/vin
+ VCTRL VCTRL VCTRL VSRC VINJ VSRC VINJ VINJ tg5v0_0[9]/vin VTUN vb VTUN VINJ VTUN
+ VTUN VINJ VINJ tg5v0_0[3]/vin l_row_en[25] vb VSRC VSRC l_row_en[22] VINJ l_row_en[21]
+ VINJ tg5v0_0[8]/vin l_row_en[24] VTUN l_row_en[27] vb VINJ VTUN l_row_en[26] VCTRL
+ VCTRL VCTRL vb VSRC tg5v0_0[2]/vin l_row_en[29] VSRC VINJ tg5v0_0[2]/vin VTUN VINJ
+ VINJ tg5v0_0[7]/vin VCTRL VCTRL VCTRL vb VTUN VSRC tg5v0_0[7]/vin VTUN vb VSRC VINJ
+ l_row_en_b[21] VINJ tg5v0_0[1]/vin l_row_en_b[28] VINJ VINJ vb VTUN l_row_en_b[25]
+ VSRC VTUN tg5v0_0[6]/vin vb VSRC VINJ VTUN l_row_en[21] VINJ VSRC l_row_en[24] l_row_en[20]
+ tg5v0_0[0]/vin l_row_en_b[25] VINJ l_row_en[23] VINJ VINJ tg5v0_0[0]/vin VCTRL VTUN
+ VINJ l_row_en[26] VCTRL VCTRL vb VSRC VTUN VSRC l_row_en[29] tg5v0_0[5]/vin vb VSRC
+ l_row_en[28] VINJ tg5v0_0[5]/vin l_row_en_b[22] VCTRL VCTRL VCTRL VTUN VINJ vb VTUN
+ VINJ VINJ l_row_en_b[29] VSRC VSRC vb VSRC VINJ l_row_en_b[22] VINJ tg5v0_0[4]/vin
+ l_row_en_b[29] VINJ VINJ VTUN l_row_en_b[26] vb VSRC VSRC tg5v0_0[9]/vin VSRC vb
+ l_row_en[20] VTUN l_row_en[23] VINJ VINJ l_row_en_b[26] tg5v0_0[3]/vin VCTRL VCTRL
+ l_row_en[22] VTUN VINJ tg5v0_0[3]/vin vb VTUN l_row_en_b[23] VSRC VSRC VINJ l_row_en[28]
+ tg5v0_0[8]/vin vb l_row_en[27] VINJ VINJ tg5v0_0[8]/vin VCTRL VCTRL VCTRL VCTRL
+ VINJ l_row_en_b[23] VINJ VINJ VTUN tg5v0_0[2]/vin l_row_en_b[24] VTUN vb VTUN VSRC
+ l_row_en_b[20] VSRC VINJ VCTRL VCTRL vb l_row_en_b[27] l_row_en_b[24] VINJ tg5v0_0[7]/vin
+ VTUN VINJ l_row_en_b[20] VINJ VINJ VINJ l_row_en_b[21] VSRC tg5v0_0[1]/vin l_row_en_b[27]
+ VTUN VSRC VSRC l_row_en[20] l_row_en_b[28] vb l_row_en_b[24] VINJ l_row_en_b[21]
+ l_row_en[22] VINJ VINJ tg5v0_0[6]/vin VTUN VINJ VTUN l_row_en_b[28] l_row_en[25]
+ vb VSRC VINJ tg5v0_0[0]/vin l_row_en[24] l_row_en_b[24] VINJ l_row_en[27] VSRC VINJ
+ tg5v0_0[0]/vin VCTRL VCTRL VCTRL VINJ VINJ l_row_en[29] tg5v0_0[5]/vin VINJ VTUN
+ l_row_en_b[25] vb VINJ tg5v0_0[5]/vin VSRC l_row_en_b[21] l_row_en[25] VCTRL VCTRL
+ VCTRL vb VSRC VSRC VINJ VTUN l_row_en_b[28] l_row_en_b[25] VTUN VINJ l_row_en_b[21]
+ VTUN VINJ VINJ VTUN VINJ l_row_en_b[22] vb VSRC l_row_en_b[28] tg5v0_0[4]/vin VSRC
+ vb l_row_en_b[29] l_row_en[22] l_row_en_b[25] vb VINJ l_row_en_b[22] l_row_en[21]
+ tg5v0_0[9]/vin VTUN VINJ l_row_en[24] VTUN VINJ l_row_en_b[29] vb l_row_en[23] tg5v0_0[3]/vin
+ l_row_en[27] VSRC l_row_en_b[25] VSRC VINJ l_row_en[26] VCTRL VCTRL VCTRL vb l_row_en_b[26]
+ VINJ VINJ l_row_en[29] tg5v0_0[3]/vin vb VTUN VINJ l_row_en_b[22] l_row_en[28] tg5v0_0[8]/vin
+ VINJ VINJ VTUN l_row_en_b[29] VSRC l_row_en_b[26] VTUN VINJ tg5v0_0[8]/vin VCTRL
+ VCTRL VCTRL vb VSRC l_row_en_b[22] vb VINJ l_row_en_b[23] tg5v0_0[2]/vin l_row_en_b[29]
+ vb VINJ VINJ VTUN VINJ l_row_en_b[26] VTUN VSRC l_row_en_b[23] vb VINJ tg5v0_0[7]/vin
+ VSRC vb tg5v0_0[1]/vin l_row_en[21] l_row_en_b[20] VINJ l_row_en_b[26] vb VINJ l_row_en[20]
+ l_row_en_b[27] VINJ tg5v0_0[1]/vin l_row_en[23] VTUN VINJ VINJ VSRC l_row_en_b[23]
+ VCTRL VCTRL VINJ l_row_en[26] l_row_en_b[20] tg5v0_0[6]/vin VCTRL vb VSRC VSRC l_row_en[25]
+ l_row_en_b[27] vb l_row_en[28] tg5v0_0[6]/vin l_row_en_b[23] VINJ vb VINJ VINJ VINJ
+ VTUN VCTRL VCTRL VINJ VINJ tg5v0_0[0]/vin VCTRL VCTRL VTUN VINJ VSRC VINJ vb VSRC
+ vb l_row_en_b[24] tg5v0_0[5]/vin l_row_en_b[20] vb VINJ VINJ VCTRL VTUN VINJ VINJ
+ VTUN l_row_en_b[27] VSRC VINJ VINJ l_row_en_b[24] VINJ vb VTUN VSRC l_row_en_b[20]
+ VINJ vb l_row_en_b[21] tg5v0_0[4]/vin l_row_en[20] l_row_en_b[27] VINJ l_row_en[23]
+ vb VTUN VINJ l_row_en_b[28] VTUN VINJ l_row_en[22] VCTRL VTUN VSRC l_row_en_b[24]
+ VINJ VSRC VINJ VINJ l_row_en_b[21] tg5v0_0[9]/vin l_row_en[25] vb VTUN l_row_en[28]
+ l_row_en_b[28] vb l_row_en[27] tg5v0_0[3]/vin l_row_en_b[24] VINJ VCTRL VCTRL VCTRL
+ vb VINJ VINJ VTUN VTUN l_row_en_b[25] VSRC VINJ VINJ tg5v0_0[3]/vin VTUN VINJ l_row_en_b[21]
+ VSRC tg5v0_0[8]/vin VINJ l_row_en_b[28] l_row_en_b[25] tg5v0_0[8]/vin VCTRL VCTRL
+ vb VINJ l_row_en_b[21] VINJ vb VTUN VINJ VTUN VSRC l_row_en_b[22] tg5v0_0[2]/vin
+ VTUN VSRC VINJ l_row_en_b[28] l_row_en[25] vb VINJ VSRC l_row_en_b[29] VINJ l_row_en[20]
+ VINJ VINJ l_row_en_b[25] VINJ l_row_en_b[22] tg5v0_0[7]/vin VINJ l_row_en[22] vb
+ VINJ VINJ l_row_en_b[29] VTUN VTUN l_row_en[25] VSRC VSRC tg5v0_0[1]/vin l_row_en_b[25]
+ l_row_en[21] VINJ vb VSRC l_row_en[24] VINJ l_row_en_b[26] tg5v0_0[1]/vin l_row_en[27]
+ l_row_en[25] vb l_row_en_b[22] l_row_en[26] VCTRL VCTRL VCTRL VINJ tg5v0_0[6]/vin
+ VINJ l_row_en[29] l_row_en_b[29] VTUN VINJ l_row_en_b[26] VTUN VSRC VINJ tg5v0_0[6]/vin
+ VSRC VINJ l_row_en_b[22] vb VTUN VSRC tg5v0_0[0]/vin VCTRL VCTRL VCTRL vb l_row_en_b[29]
+ l_row_en[25] vb VINJ VTUN VINJ VINJ VTUN VTUN l_row_en_b[23] tg5v0_0[5]/vin VSRC
+ VSRC VINJ vb VTUN VINJ VINJ l_row_en_b[26] vb VTUN VINJ l_row_en_b[23] VINJ vb VTUN
+ VINJ l_row_en[21] VINJ VTUN VINJ l_row_en[24] l_row_en_b[20] VTUN VSRC VINJ l_row_en_b[26]
+ tg5v0_0[4]/vin VSRC VINJ vb VINJ l_row_en[23] l_row_en_b[27] VINJ l_row_en[26] tg5v0_0[4]/vin
+ VCTRL VCTRL VCTRL VCTRL vb l_row_en_b[23] VINJ l_row_en[29] l_row_en_b[20] tg5v0_0[9]/vin
+ vb VINJ VTUN VSRC l_row_en[28] VSRC l_row_en_b[27] tg5v0_0[9]/vin VTUN VTUN VSRC
+ VSRC l_row_en_b[23] VCTRL VINJ VINJ VCTRL VCTRL VCTRL vb VINJ VINJ tg5v0_0[3]/vin
+ l_row_en_b[24] vb VINJ l_row_en_b[20] vb VTUN VINJ l_row_en_b[27] VSRC VSRC VTUN
+ tg5v0_0[8]/vin l_row_en_b[24] VSRC VSRC VINJ VINJ l_row_en_b[20] vb VINJ l_row_en_b[21]
+ VINJ tg5v0_0[2]/vin l_row_en_b[27] vb VINJ VGND VINJ VINJ l_row_en[21] l_row_en_b[28]
+ vb VINJ array_core_block2
Xvb_divider_0 VINJ VGND vb vb_divider
Xarray_core_block0_0 vb VINJ VTUN VTUN tg5v0_0[9]/vin VSRC l_row_en[1] VSRC VCTRL
+ l_row_en[0] tg5v0_0[3]/vin vb l_row_en[3] vb VINJ VINJ l_row_en[6] VTUN tg5v0_0[3]/vin
+ l_row_en[9] VTUN l_row_en[5] VSRC tg5v0_0[8]/vin l_row_en[8] VSRC tg5v0_0[8]/vin
+ VCTRL vb vb VINJ tg5v0_0[2]/vin VTUN VSRC VINJ VSRC VCTRL VCTRL VCTRL VINJ tg5v0_0[7]/vin
+ vb vb VINJ VTUN tg5v0_0[1]/vin VSRC VTUN VCTRL VCTRL l_row_en[0] tg5v0_0[1]/vin
+ l_row_en[3] tg5v0_0[6]/vin vb l_row_en[2] l_row_en[5] tg5v0_0[6]/vin vb VTUN VINJ
+ VINJ l_row_en[8] VSRC VSRC tg5v0_0[0]/vin l_row_en[7] vb vb VINJ tg5v0_0[5]/vin
+ VTUN VINJ VSRC VCTRL VCTRL VCTRL VCTRL VSRC VTUN vb vb tg5v0_0[4]/vin VCTRL VCTRL
+ VCTRL VCTRL l_row_en[0] VSRC VSRC l_row_en[2] tg5v0_0[9]/vin vb l_row_en[5] VTUN
+ l_row_en[4] vb tg5v0_0[3]/vin VTUN l_row_en[7] VSRC tg5v0_0[3]/vin l_row_en[9] tg5v0_0[8]/vin
+ vb VTUN tg5v0_0[8]/vin vb VTUN VCTRL VCTRL VCTRL VINJ VINJ VINJ tg5v0_0[2]/vin VCTRL
+ VCTRL VCTRL vb VSRC tg5v0_0[7]/vin VINJ VSRC l_row_en[2] tg5v0_0[1]/vin l_row_en[1]
+ vb VINJ VINJ tg5v0_0[1]/vin VTUN l_row_en[7] l_row_en[3] VSRC tg5v0_0[6]/vin VINJ
+ l_row_en[6] VSRC VINJ l_row_en[9] tg5v0_0[6]/vin l_row_en[8] vb VINJ tg5v0_0[0]/vin
+ VCTRL VCTRL vb VTUN VSRC VSRC VINJ tg5v0_0[5]/vin VCTRL VCTRL VCTRL vb VINJ VTUN
+ VINJ vb VTUN VSRC vb VINJ VINJ VINJ l_row_en[1] tg5v0_0[4]/vin VCTRL l_row_en[0]
+ vb VINJ l_row_en[3] tg5v0_0[4]/vin VTUN vb l_row_en[6] tg5v0_0[9]/vin VSRC vb VINJ
+ l_row_en[5] VINJ VINJ tg5v0_0[9]/vin l_row_en[8] VINJ VCTRL vb VINJ VTUN tg5v0_0[3]/vin
+ VSRC VINJ vb VTUN VSRC vb tg5v0_0[8]/vin VCTRL VCTRL VCTRL VCTRL VINJ VINJ vb VINJ
+ tg5v0_0[2]/vin VTUN vb VTUN VSRC VINJ vb VINJ VCTRL VCTRL VCTRL l_row_en[0] VTUN
+ tg5v0_0[7]/vin VINJ l_row_en[3] VINJ vb VINJ l_row_en[2] VTUN tg5v0_0[1]/vin VSRC
+ l_row_en[5] vb VSRC l_row_en[8] VINJ tg5v0_0[1]/vin vb VINJ l_row_en[7] VTUN tg5v0_0[6]/vin
+ VINJ vb VTUN VINJ tg5v0_0[6]/vin VTUN vb VTUN VSRC VINJ VSRC vb tg5v0_0[0]/vin VCTRL
+ VCTRL VCTRL VINJ VINJ VINJ VTUN vb VINJ VINJ tg5v0_0[5]/vin VTUN VSRC vb VCTRL VCTRL
+ VCTRL VSRC VINJ l_row_en[0] vb VINJ VINJ VTUN l_row_en[2] VINJ VINJ vb l_row_en[5]
+ l_row_en[1] VTUN VSRC tg5v0_0[4]/vin l_row_en[4] vb VSRC l_row_en[7] tg5v0_0[4]/vin
+ vb l_row_en[6] tg5v0_0[9]/vin l_row_en[9] VINJ l_row_en_b[9] VTUN VSRC VINJ tg5v0_0[9]/vin
+ VTUN VSRC l_row_en_b[2] VSRC VCTRL vb VCTRL VCTRL VTUN tg5v0_0[3]/vin VINJ VINJ
+ l_row_en_b[9] vb VINJ vb VINJ VINJ l_row_en_b[6] VTUN VSRC tg5v0_0[8]/vin VCTRL
+ VCTRL VTUN VSRC VCTRL VSRC VINJ VINJ l_row_en_b[6] tg5v0_0[2]/vin vb VINJ VINJ tg5v0_0[2]/vin
+ l_row_en[1] vb VINJ VINJ l_row_en_b[3] VTUN l_row_en[4] VTUN VSRC VSRC tg5v0_0[7]/vin
+ vb VINJ l_row_en[3] VSRC l_row_en[6] tg5v0_0[7]/vin l_row_en_b[3] l_row_en[9] VINJ
+ tg5v0_0[1]/vin l_row_en[8] vb VINJ VINJ l_row_en_b[0] VTUN VSRC VCTRL VCTRL vb VTUN
+ VSRC VINJ VSRC l_row_en_b[7] vb tg5v0_0[6]/vin VINJ VINJ l_row_en_b[0] VTUN VINJ
+ VINJ VINJ tg5v0_0[0]/vin VCTRL VCTRL VCTRL VCTRL vb l_row_en_b[7] VTUN VSRC VSRC
+ vb vb tg5v0_0[5]/vin VINJ l_row_en[1] VCTRL VCTRL VINJ VINJ l_row_en[0] vb VINJ
+ l_row_en_b[4] VINJ l_row_en[3] VTUN VTUN VSRC vb VINJ l_row_en[6] VTUN VINJ l_row_en[5]
+ vb l_row_en_b[4] tg5v0_0[4]/vin VINJ l_row_en[8] VINJ l_row_en_b[5] tg5v0_0[4]/vin
+ vb VSRC l_row_en_b[1] VTUN VINJ VSRC VSRC tg5v0_0[9]/vin vb l_row_en_b[8] l_row_en_b[5]
+ tg5v0_0[9]/vin vb VINJ l_row_en_b[1] VTUN VCTRL VCTRL VCTRL VINJ l_row_en_b[2] VTUN
+ tg5v0_0[3]/vin l_row_en_b[8] vb VSRC VINJ VINJ l_row_en_b[9] vb VSRC VINJ l_row_en_b[5]
+ l_row_en_b[2] vb tg5v0_0[8]/vin VCTRL VCTRL VCTRL l_row_en[0] VINJ VINJ l_row_en_b[9]
+ l_row_en[3] VINJ tg5v0_0[2]/vin l_row_en_b[5] vb VTUN VSRC VINJ l_row_en[2] VSRC
+ VSRC l_row_en_b[6] tg5v0_0[2]/vin l_row_en[5] vb VTUN VINJ l_row_en_b[2] l_row_en[8]
+ VTUN l_row_en[4] vb tg5v0_0[7]/vin VINJ l_row_en[7] VTUN l_row_en_b[9] l_row_en_b[6]
+ tg5v0_0[7]/vin vb VSRC l_row_en_b[2] l_row_en[9] VSRC VINJ vb tg5v0_0[1]/vin l_row_en_b[9]
+ l_row_en_b[3] VTUN VINJ vb VCTRL VCTRL VCTRL VINJ l_row_en_b[6] VTUN l_row_en_b[3]
+ VTUN tg5v0_0[6]/vin VINJ VINJ vb VSRC VTUN VINJ VSRC vb tg5v0_0[0]/vin l_row_en_b[6]
+ VCTRL VCTRL VCTRL vb VINJ tg5v0_0[0]/vin VINJ VTUN l_row_en[2] l_row_en_b[0] VSRC
+ VINJ tg5v0_0[5]/vin VSRC l_row_en[1] l_row_en[4] l_row_en_b[7] tg5v0_0[5]/vin vb
+ VINJ l_row_en[7] l_row_en_b[3] l_row_en_b[0] vb VTUN VINJ VINJ VINJ l_row_en[6]
+ VINJ VTUN l_row_en_b[7] l_row_en[9] VSRC VINJ VINJ l_row_en_b[3] VSRC VINJ l_row_en_b[4]
+ tg5v0_0[4]/vin VCTRL VCTRL l_row_en_b[0] VCTRL vb VINJ VINJ VINJ VINJ l_row_en_b[7]
+ VTUN VSRC l_row_en[4] l_row_en_b[4] VSRC tg5v0_0[9]/vin l_row_en_b[0] VSRC VCTRL
+ VCTRL vb VTUN VCTRL VCTRL VINJ l_row_en_b[1] tg5v0_0[3]/vin l_row_en_b[7] VINJ VINJ
+ l_row_en_b[8] VTUN VINJ l_row_en[1] VTUN tg5v0_0[8]/vin l_row_en_b[1] VSRC VCTRL
+ l_row_en[4] VSRC VINJ VINJ vb l_row_en[3] l_row_en_b[8] VINJ tg5v0_0[2]/vin l_row_en_b[4]
+ l_row_en[6] vb VINJ VINJ VINJ l_row_en_b[5] VTUN tg5v0_0[2]/vin l_row_en[9] VTUN
+ VINJ VTUN VINJ l_row_en_b[1] l_row_en[8] VSRC tg5v0_0[7]/vin VSRC VINJ l_row_en_b[8]
+ VCTRL vb VINJ l_row_en_b[5] VINJ tg5v0_0[7]/vin VINJ l_row_en_b[1] vb VINJ VINJ
+ VTUN VINJ l_row_en_b[2] VTUN tg5v0_0[1]/vin l_row_en_b[8] VTUN VSRC VTUN VCTRL VCTRL
+ VCTRL VSRC l_row_en_b[9] l_row_en_b[5] vb VINJ l_row_en_b[2] VTUN tg5v0_0[6]/vin
+ VINJ VINJ vb VINJ VINJ VINJ l_row_en_b[9] l_row_en[1] VTUN VTUN tg5v0_0[0]/vin VCTRL
+ VCTRL l_row_en_b[5] VTUN VSRC l_row_en[0] VSRC tg5v0_0[0]/vin l_row_en[3] vb VINJ
+ l_row_en[2] l_row_en[6] tg5v0_0[5]/vin l_row_en[5] vb VINJ VINJ VINJ VINJ l_row_en_b[6]
+ VTUN VINJ l_row_en[8] tg5v0_0[5]/vin VTUN l_row_en_b[2] VSRC VSRC VINJ VINJ l_row_en[7]
+ VTUN VTUN VSRC l_row_en_b[9] l_row_en_b[6] vb VINJ l_row_en_b[2] vb VINJ VINJ VINJ
+ VINJ l_row_en_b[3] VTUN VTUN l_row_en_b[9] tg5v0_0[4]/vin VCTRL VCTRL VCTRL VSRC
+ VSRC VINJ VSRC VINJ l_row_en_b[6] vb l_row_en_b[3] tg5v0_0[9]/vin VINJ VINJ vb VINJ
+ VINJ VCTRL VCTRL VCTRL VTUN VINJ l_row_en[0] VTUN VINJ VINJ tg5v0_0[3]/vin l_row_en_b[0]
+ VTUN l_row_en_b[6] VSRC VSRC VINJ l_row_en_b[7] VSRC VINJ l_row_en[2] tg5v0_0[3]/vin
+ VINJ l_row_en_b[3] l_row_en[5] vb tg5v0_0[8]/vin l_row_en_b[0] l_row_en[4] vb VINJ
+ VINJ VTUN l_row_en_b[7] VTUN VINJ l_row_en[7] tg5v0_0[8]/vin VTUN VTUN l_row_en_b[3]
+ VSRC VTUN VSRC l_row_en_b[4] l_row_en[9] tg5v0_0[2]/vin l_row_en_b[0] vb VINJ VINJ
+ VINJ VCTRL vb VTUN l_row_en_b[7] VCTRL VCTRL VCTRL VINJ tg5v0_0[7]/vin l_row_en_b[4]
+ VTUN VTUN VSRC l_row_en_b[0] VSRC tg5v0_0[1]/vin l_row_en_b[1] l_row_en_b[7] VSRC
+ VINJ VINJ VCTRL vb VINJ l_row_en_b[8] VCTRL VCTRL VCTRL vb VINJ VINJ VINJ VTUN l_row_en_b[4]
+ VSRC l_row_en_b[1] tg5v0_0[6]/vin VTUN VTUN l_row_en[2] VSRC VSRC l_row_en_b[8]
+ l_row_en[1] tg5v0_0[0]/vin l_row_en_b[4] VINJ l_row_en[4] VSRC VINJ VINJ VINJ l_row_en[7]
+ VINJ VINJ tg5v0_0[0]/vin vb VTUN VINJ l_row_en[6] VTUN VSRC VINJ tg5v0_0[5]/vin
+ VSRC l_row_en[9] VSRC l_row_en_b[5] tg5v0_0[5]/vin vb l_row_en_b[1] VINJ l_row_en_b[4]
+ VCTRL VCTRL VSRC VINJ VINJ VINJ l_row_en_b[8] VTUN VINJ l_row_en_b[5] VSRC VINJ
+ VTUN VINJ l_row_en_b[1] VSRC VSRC VGND VINJ l_row_en[4] l_row_en_b[2] tg5v0_0[4]/vin
+ VCTRL VCTRL vb l_row_en_b[8] VCTRL array_core_block0
.ends

.subckt top_fgcaptest vccd2 vssd2 addr[0] addr[1] addr[2] addr[3] addr[4] addr[5]
+ addr[6] addr[7] addr[8]
Xpad_minesd_short_0 VCTRL array_core_0/VCTRL array_core_0/VINJ vssd2 pad_minesd_short
Xpad_minesd_short_1 VSRC array_core_0/VSRC array_core_0/VINJ vssd2 pad_minesd_short
Xpad_minesd_short_2 VINJ array_core_0/VINJ array_core_0/VINJ vssd2 pad_minesd_short
Xpad_minesd_short_3 VOUT0 array_core_0/VOUT0 array_core_0/VINJ vssd2 pad_minesd_short
Xpad_minesd_short_4 VOUT1 array_core_0/r_vout array_core_0/VINJ vssd2 pad_minesd_short
Xvtun_pad_0 vtun_pad_0/pad vssd2 VTUN vssd2 vtun_pad
Xarray_core_0 vccd2 addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7]
+ addr[8] vtun_pad_0/pad array_core_0/VINJ array_core_0/VCTRL array_core_0/VSRC array_core_0/c[8]
+ array_core_0/c[11] array_core_0/c[14] array_core_0/c[2] array_core_0/c[7] array_core_0/c[5]
+ array_core_0/c[10] array_core_0/c[13] array_core_0/c[6] array_core_0/c[4] array_core_0/c[1]
+ array_core_0/c[9] array_core_0/r_vout array_core_0/c[12] array_core_0/VOUT0 array_core_0/c[15]
+ array_core_0/c[0] vssd2 array_core_0/c[3] array_core
.ends

