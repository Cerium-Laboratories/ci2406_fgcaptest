magic
tech sky130A
timestamp 1717562480
<< pwell >>
rect -15584 -2717 15584 2717
<< psubdiff >>
rect -15566 2682 -15518 2699
rect 15518 2682 15566 2699
rect -15566 2651 -15549 2682
rect 15549 2651 15566 2682
rect -15566 -2682 -15549 -2651
rect 15549 -2682 15566 -2651
rect -15566 -2699 -15518 -2682
rect 15518 -2699 15566 -2682
<< psubdiffcont >>
rect -15518 2682 15518 2699
rect -15566 -2651 -15549 2651
rect 15549 -2651 15566 2651
rect -15518 -2699 15518 -2682
<< xpolycontact >>
rect -15501 -2634 -14928 -2418
rect 14928 -2634 15501 -2418
<< xpolyres >>
rect -15501 2061 -14307 2634
rect -15501 -2418 -14928 2061
rect -14880 -1793 -14307 2061
rect -14259 2061 -13065 2634
rect -14259 -1793 -13686 2061
rect -14880 -2366 -13686 -1793
rect -13638 -1793 -13065 2061
rect -13017 2061 -11823 2634
rect -13017 -1793 -12444 2061
rect -13638 -2366 -12444 -1793
rect -12396 -1793 -11823 2061
rect -11775 2061 -10581 2634
rect -11775 -1793 -11202 2061
rect -12396 -2366 -11202 -1793
rect -11154 -1793 -10581 2061
rect -10533 2061 -9339 2634
rect -10533 -1793 -9960 2061
rect -11154 -2366 -9960 -1793
rect -9912 -1793 -9339 2061
rect -9291 2061 -8097 2634
rect -9291 -1793 -8718 2061
rect -9912 -2366 -8718 -1793
rect -8670 -1793 -8097 2061
rect -8049 2061 -6855 2634
rect -8049 -1793 -7476 2061
rect -8670 -2366 -7476 -1793
rect -7428 -1793 -6855 2061
rect -6807 2061 -5613 2634
rect -6807 -1793 -6234 2061
rect -7428 -2366 -6234 -1793
rect -6186 -1793 -5613 2061
rect -5565 2061 -4371 2634
rect -5565 -1793 -4992 2061
rect -6186 -2366 -4992 -1793
rect -4944 -1793 -4371 2061
rect -4323 2061 -3129 2634
rect -4323 -1793 -3750 2061
rect -4944 -2366 -3750 -1793
rect -3702 -1793 -3129 2061
rect -3081 2061 -1887 2634
rect -3081 -1793 -2508 2061
rect -3702 -2366 -2508 -1793
rect -2460 -1793 -1887 2061
rect -1839 2061 -645 2634
rect -1839 -1793 -1266 2061
rect -2460 -2366 -1266 -1793
rect -1218 -1793 -645 2061
rect -597 2061 597 2634
rect -597 -1793 -24 2061
rect -1218 -2366 -24 -1793
rect 24 -1793 597 2061
rect 645 2061 1839 2634
rect 645 -1793 1218 2061
rect 24 -2366 1218 -1793
rect 1266 -1793 1839 2061
rect 1887 2061 3081 2634
rect 1887 -1793 2460 2061
rect 1266 -2366 2460 -1793
rect 2508 -1793 3081 2061
rect 3129 2061 4323 2634
rect 3129 -1793 3702 2061
rect 2508 -2366 3702 -1793
rect 3750 -1793 4323 2061
rect 4371 2061 5565 2634
rect 4371 -1793 4944 2061
rect 3750 -2366 4944 -1793
rect 4992 -1793 5565 2061
rect 5613 2061 6807 2634
rect 5613 -1793 6186 2061
rect 4992 -2366 6186 -1793
rect 6234 -1793 6807 2061
rect 6855 2061 8049 2634
rect 6855 -1793 7428 2061
rect 6234 -2366 7428 -1793
rect 7476 -1793 8049 2061
rect 8097 2061 9291 2634
rect 8097 -1793 8670 2061
rect 7476 -2366 8670 -1793
rect 8718 -1793 9291 2061
rect 9339 2061 10533 2634
rect 9339 -1793 9912 2061
rect 8718 -2366 9912 -1793
rect 9960 -1793 10533 2061
rect 10581 2061 11775 2634
rect 10581 -1793 11154 2061
rect 9960 -2366 11154 -1793
rect 11202 -1793 11775 2061
rect 11823 2061 13017 2634
rect 11823 -1793 12396 2061
rect 11202 -2366 12396 -1793
rect 12444 -1793 13017 2061
rect 13065 2061 14259 2634
rect 13065 -1793 13638 2061
rect 12444 -2366 13638 -1793
rect 13686 -1793 14259 2061
rect 14307 2061 15501 2634
rect 14307 -1793 14880 2061
rect 13686 -2366 14880 -1793
rect 14928 -2418 15501 2061
<< locali >>
rect -15566 2682 -15518 2699
rect 15518 2682 15566 2699
rect -15566 2651 -15549 2682
rect 15549 2651 15566 2682
rect -15566 -2682 -15549 -2651
rect 15549 -2682 15566 -2651
rect -15566 -2699 -15518 -2682
rect 15518 -2699 15566 -2682
<< properties >>
string FIXED_BBOX -15557 -2690 15557 2690
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 50 m 1 nx 50 wmin 5.730 lmin 0.50 rho 2000 val 970.666k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
