magic
tech sky130A
timestamp 1717158785
<< error_p >>
rect 349 13678 580 13758
rect 2349 13678 2580 13758
rect 4349 13678 4580 13758
rect 6349 13678 6580 13758
rect 8349 13678 8580 13758
rect 10349 13678 10580 13758
rect 12349 13678 12580 13758
rect 14349 13678 14580 13758
rect 16349 13678 16580 13758
rect 18349 13678 18580 13758
rect 349 12178 580 12258
rect 2349 12178 2580 12258
rect 4349 12178 4580 12258
rect 6349 12178 6580 12258
rect 8349 12178 8580 12258
rect 10349 12178 10580 12258
rect 12349 12178 12580 12258
rect 14349 12178 14580 12258
rect 16349 12178 16580 12258
rect 18349 12178 18580 12258
rect 349 10678 580 10758
rect 2349 10678 2580 10758
rect 4349 10678 4580 10758
rect 6349 10678 6580 10758
rect 8349 10678 8580 10758
rect 10349 10678 10580 10758
rect 12349 10678 12580 10758
rect 14349 10678 14580 10758
rect 16349 10678 16580 10758
rect 18349 10678 18580 10758
rect 349 9178 580 9258
rect 2349 9178 2580 9258
rect 4349 9178 4580 9258
rect 6349 9178 6580 9258
rect 8349 9178 8580 9258
rect 10349 9178 10580 9258
rect 12349 9178 12580 9258
rect 14349 9178 14580 9258
rect 16349 9178 16580 9258
rect 18349 9178 18580 9258
rect 349 7678 580 7758
rect 2349 7678 2580 7758
rect 4349 7678 4580 7758
rect 6349 7678 6580 7758
rect 8349 7678 8580 7758
rect 10349 7678 10580 7758
rect 12349 7678 12580 7758
rect 14349 7678 14580 7758
rect 16349 7678 16580 7758
rect 18349 7678 18580 7758
rect 349 6178 580 6258
rect 2349 6178 2580 6258
rect 4349 6178 4580 6258
rect 6349 6178 6580 6258
rect 8349 6178 8580 6258
rect 10349 6178 10580 6258
rect 12349 6178 12580 6258
rect 14349 6178 14580 6258
rect 16349 6178 16580 6258
rect 18349 6178 18580 6258
rect 349 4678 580 4758
rect 2349 4678 2580 4758
rect 4349 4678 4580 4758
rect 6349 4678 6580 4758
rect 8349 4678 8580 4758
rect 10349 4678 10580 4758
rect 12349 4678 12580 4758
rect 14349 4678 14580 4758
rect 16349 4678 16580 4758
rect 18349 4678 18580 4758
rect 349 3178 580 3258
rect 2349 3178 2580 3258
rect 4349 3178 4580 3258
rect 6349 3178 6580 3258
rect 8349 3178 8580 3258
rect 10349 3178 10580 3258
rect 12349 3178 12580 3258
rect 14349 3178 14580 3258
rect 16349 3178 16580 3258
rect 18349 3178 18580 3258
rect 349 1678 580 1758
rect 2349 1678 2580 1758
rect 4349 1678 4580 1758
rect 6349 1678 6580 1758
rect 8349 1678 8580 1758
rect 10349 1678 10580 1758
rect 12349 1678 12580 1758
rect 14349 1678 14580 1758
rect 16349 1678 16580 1758
rect 18349 1678 18580 1758
rect 349 178 580 258
rect 2349 178 2580 258
rect 4349 178 4580 258
rect 6349 178 6580 258
rect 8349 178 8580 258
rect 10349 178 10580 258
rect 12349 178 12580 258
rect 14349 178 14580 258
rect 16349 178 16580 258
rect 18349 178 18580 258
use fgcell_amp_MiM_cap_1_1  fgcell_amp_MiM_cap_1_1_0
array 0 9 2000 0 9 1500
timestamp 1717158785
transform 1 0 -262 0 1 1403
box 262 -2099 2245 -785
<< end >>
