magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< pwell >>
rect 0 0 1518 1972
<< mvpsubdiff >>
rect 66 1894 1452 1906
rect 66 1860 174 1894
rect 1368 1860 1452 1894
rect 66 1848 1452 1860
rect 66 1798 124 1848
rect 66 174 78 1798
rect 112 174 124 1798
rect 1394 1798 1452 1848
rect 66 124 124 174
rect 1394 174 1406 1798
rect 1440 174 1452 1798
rect 1394 124 1452 174
rect 66 112 1452 124
rect 66 78 174 112
rect 1368 78 1452 112
rect 66 66 1452 78
<< mvpsubdiffcont >>
rect 174 1860 1368 1894
rect 78 174 112 1798
rect 1406 174 1440 1798
rect 174 78 1368 112
<< xpolycontact >>
rect 220 1320 290 1752
rect 220 220 290 652
rect 332 1320 402 1752
rect 332 220 402 652
rect 444 1320 514 1752
rect 444 220 514 652
rect 556 1320 626 1752
rect 556 220 626 652
rect 668 1320 738 1752
rect 668 220 738 652
rect 780 1320 850 1752
rect 780 220 850 652
rect 892 1320 962 1752
rect 892 220 962 652
rect 1004 1320 1074 1752
rect 1004 220 1074 652
rect 1116 1320 1186 1752
rect 1116 220 1186 652
rect 1228 1320 1298 1752
rect 1228 220 1298 652
<< xpolyres >>
rect 220 652 290 1320
rect 332 652 402 1320
rect 444 652 514 1320
rect 556 652 626 1320
rect 668 652 738 1320
rect 780 652 850 1320
rect 892 652 962 1320
rect 1004 652 1074 1320
rect 1116 652 1186 1320
rect 1228 652 1298 1320
<< locali >>
rect 78 1860 174 1894
rect 1368 1860 1440 1894
rect 78 1798 112 1860
rect 444 1752 514 1860
rect 1406 1798 1440 1860
rect 78 112 112 174
rect 1406 112 1440 174
rect 78 78 174 112
rect 1368 78 1440 112
<< viali >>
rect 174 1860 1368 1894
rect 236 1337 274 1734
rect 348 1337 386 1734
rect 460 1337 498 1734
rect 572 1337 610 1734
rect 684 1337 722 1734
rect 796 1337 834 1734
rect 908 1337 946 1734
rect 1020 1337 1058 1734
rect 1132 1337 1170 1734
rect 1244 1337 1282 1734
rect 236 238 274 635
rect 348 238 386 635
rect 460 238 498 635
rect 572 238 610 635
rect 684 238 722 635
rect 796 238 834 635
rect 908 238 946 635
rect 1020 238 1058 635
rect 1132 238 1170 635
rect 1244 238 1282 635
<< metal1 >>
rect 66 1894 1452 1906
rect 66 1860 174 1894
rect 1368 1860 1452 1894
rect 66 1854 1452 1860
rect 66 118 118 1854
rect 342 1776 616 1826
rect 230 1734 280 1746
rect 230 1337 236 1734
rect 274 1337 280 1734
rect 230 1325 280 1337
rect 342 1734 392 1776
rect 342 1337 348 1734
rect 386 1337 392 1734
rect 342 1324 392 1337
rect 454 1734 504 1746
rect 454 1337 460 1734
rect 498 1337 504 1734
rect 454 1324 504 1337
rect 566 1734 616 1776
rect 902 1776 1176 1826
rect 566 1337 572 1734
rect 610 1337 616 1734
rect 566 1324 616 1337
rect 678 1734 840 1746
rect 678 1337 684 1734
rect 722 1337 796 1734
rect 834 1337 840 1734
rect 678 1324 840 1337
rect 902 1734 952 1776
rect 902 1337 908 1734
rect 946 1337 952 1734
rect 902 1324 952 1337
rect 1014 1734 1064 1746
rect 1014 1337 1020 1734
rect 1058 1337 1064 1734
rect 1014 1294 1064 1337
rect 1126 1734 1176 1776
rect 1126 1337 1132 1734
rect 1170 1337 1176 1734
rect 1126 1324 1176 1337
rect 1238 1734 1288 1746
rect 1238 1337 1244 1734
rect 1282 1337 1288 1734
rect 1238 1294 1288 1337
rect 1014 1244 1288 1294
rect 230 635 392 648
rect 230 238 236 635
rect 274 238 348 635
rect 386 238 392 635
rect 230 226 392 238
rect 454 635 504 648
rect 454 238 460 635
rect 498 238 504 635
rect 454 196 504 238
rect 566 635 728 648
rect 566 238 572 635
rect 610 238 684 635
rect 722 238 728 635
rect 566 226 728 238
rect 790 635 952 648
rect 790 238 796 635
rect 834 238 908 635
rect 946 238 952 635
rect 790 226 952 238
rect 1014 635 1064 648
rect 1014 238 1020 635
rect 1058 238 1064 635
rect 1014 196 1064 238
rect 1126 635 1288 648
rect 1126 238 1132 635
rect 1170 238 1244 635
rect 1282 238 1288 635
rect 1126 226 1288 238
rect 454 146 1064 196
rect 1400 118 1452 1854
rect 66 66 1452 118
<< labels >>
flabel metal1 230 1325 280 1746 0 FreeSans 320 90 0 0 VDD
port 1 nsew power default
flabel metal1 1238 1326 1288 1746 0 FreeSans 320 90 0 0 vout_1v
port 3 nsew analog default
flabel metal1 454 1324 504 1746 0 FreeSans 320 90 0 0 VGND
port 2 nsew ground default
flabel pwell 124 1798 174 1848 0 FreeSans 160 0 0 0 VGND
flabel metal1 66 1854 118 1906 0 FreeSans 160 0 0 0 VGND
<< end >>
