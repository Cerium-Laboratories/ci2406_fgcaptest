magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< error_p >>
rect 1982 29160 2302 29230
rect 366 28916 606 28940
rect 366 28724 390 28916
rect 582 28724 606 28916
rect 1982 28920 2006 29160
rect 2232 28920 2246 29160
rect 2256 28920 2302 29160
rect 5982 29160 6302 29230
rect 1982 28896 2302 28920
rect 4366 28916 4606 28940
rect 366 28700 606 28724
rect 4366 28724 4390 28916
rect 4582 28724 4606 28916
rect 5982 28920 6006 29160
rect 6232 28920 6246 29160
rect 6256 28920 6302 29160
rect 9982 29160 10302 29230
rect 5982 28896 6302 28920
rect 8366 28916 8606 28940
rect 2852 28709 2996 28714
rect 2852 28639 2857 28709
rect 2991 28639 2996 28709
rect 4366 28700 4606 28724
rect 8366 28724 8390 28916
rect 8582 28724 8606 28916
rect 9982 28920 10006 29160
rect 10232 28920 10246 29160
rect 10256 28920 10302 29160
rect 13982 29160 14302 29230
rect 9982 28896 10302 28920
rect 12366 28916 12606 28940
rect 6852 28709 6996 28714
rect 2852 28634 2996 28639
rect 6852 28639 6857 28709
rect 6991 28639 6996 28709
rect 8366 28700 8606 28724
rect 12366 28724 12390 28916
rect 12582 28724 12606 28916
rect 13982 28920 14006 29160
rect 14232 28920 14246 29160
rect 14256 28920 14302 29160
rect 17982 29160 18302 29230
rect 13982 28896 14302 28920
rect 16366 28916 16606 28940
rect 10852 28709 10996 28714
rect 6852 28634 6996 28639
rect 10852 28639 10857 28709
rect 10991 28639 10996 28709
rect 12366 28700 12606 28724
rect 16366 28724 16390 28916
rect 16582 28724 16606 28916
rect 17982 28920 18006 29160
rect 18232 28920 18246 29160
rect 18256 28920 18302 29160
rect 21982 29160 22302 29230
rect 17982 28896 18302 28920
rect 20366 28916 20606 28940
rect 14852 28709 14996 28714
rect 10852 28634 10996 28639
rect 14852 28639 14857 28709
rect 14991 28639 14996 28709
rect 16366 28700 16606 28724
rect 20366 28724 20390 28916
rect 20582 28724 20606 28916
rect 21982 28920 22006 29160
rect 22232 28920 22246 29160
rect 22256 28920 22302 29160
rect 25982 29160 26302 29230
rect 21982 28896 22302 28920
rect 24366 28916 24606 28940
rect 18852 28709 18996 28714
rect 14852 28634 14996 28639
rect 18852 28639 18857 28709
rect 18991 28639 18996 28709
rect 20366 28700 20606 28724
rect 24366 28724 24390 28916
rect 24582 28724 24606 28916
rect 25982 28920 26006 29160
rect 26232 28920 26246 29160
rect 26256 28920 26302 29160
rect 29982 29160 30302 29230
rect 25982 28896 26302 28920
rect 28366 28916 28606 28940
rect 22852 28709 22996 28714
rect 18852 28634 18996 28639
rect 22852 28639 22857 28709
rect 22991 28639 22996 28709
rect 24366 28700 24606 28724
rect 28366 28724 28390 28916
rect 28582 28724 28606 28916
rect 29982 28920 30006 29160
rect 30232 28920 30246 29160
rect 30256 28920 30302 29160
rect 33982 29160 34302 29230
rect 29982 28896 30302 28920
rect 32366 28916 32606 28940
rect 26852 28709 26996 28714
rect 22852 28634 22996 28639
rect 26852 28639 26857 28709
rect 26991 28639 26996 28709
rect 28366 28700 28606 28724
rect 32366 28724 32390 28916
rect 32582 28724 32606 28916
rect 33982 28920 34006 29160
rect 34232 28920 34246 29160
rect 34256 28920 34302 29160
rect 37982 29160 38302 29230
rect 33982 28896 34302 28920
rect 36366 28916 36606 28940
rect 30852 28709 30996 28714
rect 26852 28634 26996 28639
rect 30852 28639 30857 28709
rect 30991 28639 30996 28709
rect 32366 28700 32606 28724
rect 36366 28724 36390 28916
rect 36582 28724 36606 28916
rect 37982 28920 38006 29160
rect 38232 28920 38246 29160
rect 38256 28920 38302 29160
rect 37982 28896 38302 28920
rect 34852 28709 34996 28714
rect 30852 28634 30996 28639
rect 34852 28639 34857 28709
rect 34991 28639 34996 28709
rect 36366 28700 36606 28724
rect 38852 28709 38996 28714
rect 34852 28634 34996 28639
rect 38852 28639 38857 28709
rect 38991 28639 38996 28709
rect 38852 28634 38996 28639
rect 2366 28559 2546 28560
rect 2366 28381 2367 28559
rect 2545 28381 2546 28559
rect 2366 28380 2546 28381
rect 6366 28559 6546 28560
rect 6366 28381 6367 28559
rect 6545 28381 6546 28559
rect 6366 28380 6546 28381
rect 10366 28559 10546 28560
rect 10366 28381 10367 28559
rect 10545 28381 10546 28559
rect 10366 28380 10546 28381
rect 14366 28559 14546 28560
rect 14366 28381 14367 28559
rect 14545 28381 14546 28559
rect 14366 28380 14546 28381
rect 18366 28559 18546 28560
rect 18366 28381 18367 28559
rect 18545 28381 18546 28559
rect 18366 28380 18546 28381
rect 22366 28559 22546 28560
rect 22366 28381 22367 28559
rect 22545 28381 22546 28559
rect 22366 28380 22546 28381
rect 26366 28559 26546 28560
rect 26366 28381 26367 28559
rect 26545 28381 26546 28559
rect 26366 28380 26546 28381
rect 30366 28559 30546 28560
rect 30366 28381 30367 28559
rect 30545 28381 30546 28559
rect 30366 28380 30546 28381
rect 34366 28559 34546 28560
rect 34366 28381 34367 28559
rect 34545 28381 34546 28559
rect 34366 28380 34546 28381
rect 38366 28559 38546 28560
rect 38366 28381 38367 28559
rect 38545 28381 38546 28559
rect 38366 28380 38546 28381
rect 366 28039 546 28040
rect 366 27861 367 28039
rect 545 27861 546 28039
rect 4366 28039 4546 28040
rect 3734 27984 3740 27990
rect 3780 27984 3786 27990
rect 3728 27978 3734 27984
rect 3786 27978 3792 27984
rect 3728 27928 3734 27934
rect 3786 27928 3792 27934
rect 3734 27922 3740 27928
rect 3780 27922 3786 27928
rect 366 27860 546 27861
rect 4366 27861 4367 28039
rect 4545 27861 4546 28039
rect 8366 28039 8546 28040
rect 7734 27984 7740 27990
rect 7780 27984 7786 27990
rect 7728 27978 7734 27984
rect 7786 27978 7792 27984
rect 7728 27928 7734 27934
rect 7786 27928 7792 27934
rect 7734 27922 7740 27928
rect 7780 27922 7786 27928
rect 4366 27860 4546 27861
rect 8366 27861 8367 28039
rect 8545 27861 8546 28039
rect 12366 28039 12546 28040
rect 11734 27984 11740 27990
rect 11780 27984 11786 27990
rect 11728 27978 11734 27984
rect 11786 27978 11792 27984
rect 11728 27928 11734 27934
rect 11786 27928 11792 27934
rect 11734 27922 11740 27928
rect 11780 27922 11786 27928
rect 8366 27860 8546 27861
rect 12366 27861 12367 28039
rect 12545 27861 12546 28039
rect 16366 28039 16546 28040
rect 15734 27984 15740 27990
rect 15780 27984 15786 27990
rect 15728 27978 15734 27984
rect 15786 27978 15792 27984
rect 15728 27928 15734 27934
rect 15786 27928 15792 27934
rect 15734 27922 15740 27928
rect 15780 27922 15786 27928
rect 12366 27860 12546 27861
rect 16366 27861 16367 28039
rect 16545 27861 16546 28039
rect 20366 28039 20546 28040
rect 19734 27984 19740 27990
rect 19780 27984 19786 27990
rect 19728 27978 19734 27984
rect 19786 27978 19792 27984
rect 19728 27928 19734 27934
rect 19786 27928 19792 27934
rect 19734 27922 19740 27928
rect 19780 27922 19786 27928
rect 16366 27860 16546 27861
rect 20366 27861 20367 28039
rect 20545 27861 20546 28039
rect 24366 28039 24546 28040
rect 23734 27984 23740 27990
rect 23780 27984 23786 27990
rect 23728 27978 23734 27984
rect 23786 27978 23792 27984
rect 23728 27928 23734 27934
rect 23786 27928 23792 27934
rect 23734 27922 23740 27928
rect 23780 27922 23786 27928
rect 20366 27860 20546 27861
rect 24366 27861 24367 28039
rect 24545 27861 24546 28039
rect 28366 28039 28546 28040
rect 27734 27984 27740 27990
rect 27780 27984 27786 27990
rect 27728 27978 27734 27984
rect 27786 27978 27792 27984
rect 27728 27928 27734 27934
rect 27786 27928 27792 27934
rect 27734 27922 27740 27928
rect 27780 27922 27786 27928
rect 24366 27860 24546 27861
rect 28366 27861 28367 28039
rect 28545 27861 28546 28039
rect 32366 28039 32546 28040
rect 31734 27984 31740 27990
rect 31780 27984 31786 27990
rect 31728 27978 31734 27984
rect 31786 27978 31792 27984
rect 31728 27928 31734 27934
rect 31786 27928 31792 27934
rect 31734 27922 31740 27928
rect 31780 27922 31786 27928
rect 28366 27860 28546 27861
rect 32366 27861 32367 28039
rect 32545 27861 32546 28039
rect 36366 28039 36546 28040
rect 35734 27984 35740 27990
rect 35780 27984 35786 27990
rect 35728 27978 35734 27984
rect 35786 27978 35792 27984
rect 35728 27928 35734 27934
rect 35786 27928 35792 27934
rect 35734 27922 35740 27928
rect 35780 27922 35786 27928
rect 32366 27860 32546 27861
rect 36366 27861 36367 28039
rect 36545 27861 36546 28039
rect 39734 27984 39740 27990
rect 39780 27984 39786 27990
rect 39728 27978 39734 27984
rect 39786 27978 39792 27984
rect 39728 27928 39734 27934
rect 39786 27928 39792 27934
rect 39734 27922 39740 27928
rect 39780 27922 39786 27928
rect 36366 27860 36546 27861
rect 3262 27808 3268 27814
rect 3308 27808 3314 27814
rect 7262 27808 7268 27814
rect 7308 27808 7314 27814
rect 11262 27808 11268 27814
rect 11308 27808 11314 27814
rect 15262 27808 15268 27814
rect 15308 27808 15314 27814
rect 19262 27808 19268 27814
rect 19308 27808 19314 27814
rect 23262 27808 23268 27814
rect 23308 27808 23314 27814
rect 27262 27808 27268 27814
rect 27308 27808 27314 27814
rect 31262 27808 31268 27814
rect 31308 27808 31314 27814
rect 35262 27808 35268 27814
rect 35308 27808 35314 27814
rect 39262 27808 39268 27814
rect 39308 27808 39314 27814
rect 3256 27802 3262 27808
rect 3314 27802 3320 27808
rect 7256 27802 7262 27808
rect 7314 27802 7320 27808
rect 11256 27802 11262 27808
rect 11314 27802 11320 27808
rect 15256 27802 15262 27808
rect 15314 27802 15320 27808
rect 19256 27802 19262 27808
rect 19314 27802 19320 27808
rect 23256 27802 23262 27808
rect 23314 27802 23320 27808
rect 27256 27802 27262 27808
rect 27314 27802 27320 27808
rect 31256 27802 31262 27808
rect 31314 27802 31320 27808
rect 35256 27802 35262 27808
rect 35314 27802 35320 27808
rect 39256 27802 39262 27808
rect 39314 27802 39320 27808
rect 3256 27756 3262 27762
rect 3314 27756 3320 27762
rect 7256 27756 7262 27762
rect 7314 27756 7320 27762
rect 11256 27756 11262 27762
rect 11314 27756 11320 27762
rect 15256 27756 15262 27762
rect 15314 27756 15320 27762
rect 19256 27756 19262 27762
rect 19314 27756 19320 27762
rect 23256 27756 23262 27762
rect 23314 27756 23320 27762
rect 27256 27756 27262 27762
rect 27314 27756 27320 27762
rect 31256 27756 31262 27762
rect 31314 27756 31320 27762
rect 35256 27756 35262 27762
rect 35314 27756 35320 27762
rect 39256 27756 39262 27762
rect 39314 27756 39320 27762
rect 3262 27750 3268 27756
rect 3308 27750 3314 27756
rect 7262 27750 7268 27756
rect 7308 27750 7314 27756
rect 11262 27750 11268 27756
rect 11308 27750 11314 27756
rect 15262 27750 15268 27756
rect 15308 27750 15314 27756
rect 19262 27750 19268 27756
rect 19308 27750 19314 27756
rect 23262 27750 23268 27756
rect 23308 27750 23314 27756
rect 27262 27750 27268 27756
rect 27308 27750 27314 27756
rect 31262 27750 31268 27756
rect 31308 27750 31314 27756
rect 35262 27750 35268 27756
rect 35308 27750 35314 27756
rect 39262 27750 39268 27756
rect 39308 27750 39314 27756
rect 2386 27296 2626 27320
rect 2386 27104 2410 27296
rect 2602 27104 2626 27296
rect 2386 27080 2626 27104
rect 6386 27296 6626 27320
rect 6386 27104 6410 27296
rect 6602 27104 6626 27296
rect 6386 27080 6626 27104
rect 10386 27296 10626 27320
rect 10386 27104 10410 27296
rect 10602 27104 10626 27296
rect 10386 27080 10626 27104
rect 14386 27296 14626 27320
rect 14386 27104 14410 27296
rect 14602 27104 14626 27296
rect 14386 27080 14626 27104
rect 18386 27296 18626 27320
rect 18386 27104 18410 27296
rect 18602 27104 18626 27296
rect 18386 27080 18626 27104
rect 22386 27296 22626 27320
rect 22386 27104 22410 27296
rect 22602 27104 22626 27296
rect 22386 27080 22626 27104
rect 26386 27296 26626 27320
rect 26386 27104 26410 27296
rect 26602 27104 26626 27296
rect 26386 27080 26626 27104
rect 30386 27296 30626 27320
rect 30386 27104 30410 27296
rect 30602 27104 30626 27296
rect 30386 27080 30626 27104
rect 34386 27296 34626 27320
rect 34386 27104 34410 27296
rect 34602 27104 34626 27296
rect 34386 27080 34626 27104
rect 38386 27296 38626 27320
rect 38386 27104 38410 27296
rect 38602 27104 38626 27296
rect 38386 27080 38626 27104
rect 1982 26160 2302 26230
rect 366 25916 606 25940
rect 366 25724 390 25916
rect 582 25724 606 25916
rect 1982 25920 2006 26160
rect 2232 25920 2246 26160
rect 2256 25920 2302 26160
rect 5982 26160 6302 26230
rect 1982 25896 2302 25920
rect 4366 25916 4606 25940
rect 366 25700 606 25724
rect 4366 25724 4390 25916
rect 4582 25724 4606 25916
rect 5982 25920 6006 26160
rect 6232 25920 6246 26160
rect 6256 25920 6302 26160
rect 9982 26160 10302 26230
rect 5982 25896 6302 25920
rect 8366 25916 8606 25940
rect 2852 25709 2996 25714
rect 2852 25639 2857 25709
rect 2991 25639 2996 25709
rect 4366 25700 4606 25724
rect 8366 25724 8390 25916
rect 8582 25724 8606 25916
rect 9982 25920 10006 26160
rect 10232 25920 10246 26160
rect 10256 25920 10302 26160
rect 13982 26160 14302 26230
rect 9982 25896 10302 25920
rect 12366 25916 12606 25940
rect 6852 25709 6996 25714
rect 2852 25634 2996 25639
rect 6852 25639 6857 25709
rect 6991 25639 6996 25709
rect 8366 25700 8606 25724
rect 12366 25724 12390 25916
rect 12582 25724 12606 25916
rect 13982 25920 14006 26160
rect 14232 25920 14246 26160
rect 14256 25920 14302 26160
rect 17982 26160 18302 26230
rect 13982 25896 14302 25920
rect 16366 25916 16606 25940
rect 10852 25709 10996 25714
rect 6852 25634 6996 25639
rect 10852 25639 10857 25709
rect 10991 25639 10996 25709
rect 12366 25700 12606 25724
rect 16366 25724 16390 25916
rect 16582 25724 16606 25916
rect 17982 25920 18006 26160
rect 18232 25920 18246 26160
rect 18256 25920 18302 26160
rect 21982 26160 22302 26230
rect 17982 25896 18302 25920
rect 20366 25916 20606 25940
rect 14852 25709 14996 25714
rect 10852 25634 10996 25639
rect 14852 25639 14857 25709
rect 14991 25639 14996 25709
rect 16366 25700 16606 25724
rect 20366 25724 20390 25916
rect 20582 25724 20606 25916
rect 21982 25920 22006 26160
rect 22232 25920 22246 26160
rect 22256 25920 22302 26160
rect 25982 26160 26302 26230
rect 21982 25896 22302 25920
rect 24366 25916 24606 25940
rect 18852 25709 18996 25714
rect 14852 25634 14996 25639
rect 18852 25639 18857 25709
rect 18991 25639 18996 25709
rect 20366 25700 20606 25724
rect 24366 25724 24390 25916
rect 24582 25724 24606 25916
rect 25982 25920 26006 26160
rect 26232 25920 26246 26160
rect 26256 25920 26302 26160
rect 29982 26160 30302 26230
rect 25982 25896 26302 25920
rect 28366 25916 28606 25940
rect 22852 25709 22996 25714
rect 18852 25634 18996 25639
rect 22852 25639 22857 25709
rect 22991 25639 22996 25709
rect 24366 25700 24606 25724
rect 28366 25724 28390 25916
rect 28582 25724 28606 25916
rect 29982 25920 30006 26160
rect 30232 25920 30246 26160
rect 30256 25920 30302 26160
rect 33982 26160 34302 26230
rect 29982 25896 30302 25920
rect 32366 25916 32606 25940
rect 26852 25709 26996 25714
rect 22852 25634 22996 25639
rect 26852 25639 26857 25709
rect 26991 25639 26996 25709
rect 28366 25700 28606 25724
rect 32366 25724 32390 25916
rect 32582 25724 32606 25916
rect 33982 25920 34006 26160
rect 34232 25920 34246 26160
rect 34256 25920 34302 26160
rect 37982 26160 38302 26230
rect 33982 25896 34302 25920
rect 36366 25916 36606 25940
rect 30852 25709 30996 25714
rect 26852 25634 26996 25639
rect 30852 25639 30857 25709
rect 30991 25639 30996 25709
rect 32366 25700 32606 25724
rect 36366 25724 36390 25916
rect 36582 25724 36606 25916
rect 37982 25920 38006 26160
rect 38232 25920 38246 26160
rect 38256 25920 38302 26160
rect 37982 25896 38302 25920
rect 34852 25709 34996 25714
rect 30852 25634 30996 25639
rect 34852 25639 34857 25709
rect 34991 25639 34996 25709
rect 36366 25700 36606 25724
rect 38852 25709 38996 25714
rect 34852 25634 34996 25639
rect 38852 25639 38857 25709
rect 38991 25639 38996 25709
rect 38852 25634 38996 25639
rect 2366 25559 2546 25560
rect 2366 25381 2367 25559
rect 2545 25381 2546 25559
rect 2366 25380 2546 25381
rect 6366 25559 6546 25560
rect 6366 25381 6367 25559
rect 6545 25381 6546 25559
rect 6366 25380 6546 25381
rect 10366 25559 10546 25560
rect 10366 25381 10367 25559
rect 10545 25381 10546 25559
rect 10366 25380 10546 25381
rect 14366 25559 14546 25560
rect 14366 25381 14367 25559
rect 14545 25381 14546 25559
rect 14366 25380 14546 25381
rect 18366 25559 18546 25560
rect 18366 25381 18367 25559
rect 18545 25381 18546 25559
rect 18366 25380 18546 25381
rect 22366 25559 22546 25560
rect 22366 25381 22367 25559
rect 22545 25381 22546 25559
rect 22366 25380 22546 25381
rect 26366 25559 26546 25560
rect 26366 25381 26367 25559
rect 26545 25381 26546 25559
rect 26366 25380 26546 25381
rect 30366 25559 30546 25560
rect 30366 25381 30367 25559
rect 30545 25381 30546 25559
rect 30366 25380 30546 25381
rect 34366 25559 34546 25560
rect 34366 25381 34367 25559
rect 34545 25381 34546 25559
rect 34366 25380 34546 25381
rect 38366 25559 38546 25560
rect 38366 25381 38367 25559
rect 38545 25381 38546 25559
rect 38366 25380 38546 25381
rect 366 25039 546 25040
rect 366 24861 367 25039
rect 545 24861 546 25039
rect 4366 25039 4546 25040
rect 3734 24984 3740 24990
rect 3780 24984 3786 24990
rect 3728 24978 3734 24984
rect 3786 24978 3792 24984
rect 3728 24928 3734 24934
rect 3786 24928 3792 24934
rect 3734 24922 3740 24928
rect 3780 24922 3786 24928
rect 366 24860 546 24861
rect 4366 24861 4367 25039
rect 4545 24861 4546 25039
rect 8366 25039 8546 25040
rect 7734 24984 7740 24990
rect 7780 24984 7786 24990
rect 7728 24978 7734 24984
rect 7786 24978 7792 24984
rect 7728 24928 7734 24934
rect 7786 24928 7792 24934
rect 7734 24922 7740 24928
rect 7780 24922 7786 24928
rect 4366 24860 4546 24861
rect 8366 24861 8367 25039
rect 8545 24861 8546 25039
rect 12366 25039 12546 25040
rect 11734 24984 11740 24990
rect 11780 24984 11786 24990
rect 11728 24978 11734 24984
rect 11786 24978 11792 24984
rect 11728 24928 11734 24934
rect 11786 24928 11792 24934
rect 11734 24922 11740 24928
rect 11780 24922 11786 24928
rect 8366 24860 8546 24861
rect 12366 24861 12367 25039
rect 12545 24861 12546 25039
rect 16366 25039 16546 25040
rect 15734 24984 15740 24990
rect 15780 24984 15786 24990
rect 15728 24978 15734 24984
rect 15786 24978 15792 24984
rect 15728 24928 15734 24934
rect 15786 24928 15792 24934
rect 15734 24922 15740 24928
rect 15780 24922 15786 24928
rect 12366 24860 12546 24861
rect 16366 24861 16367 25039
rect 16545 24861 16546 25039
rect 20366 25039 20546 25040
rect 19734 24984 19740 24990
rect 19780 24984 19786 24990
rect 19728 24978 19734 24984
rect 19786 24978 19792 24984
rect 19728 24928 19734 24934
rect 19786 24928 19792 24934
rect 19734 24922 19740 24928
rect 19780 24922 19786 24928
rect 16366 24860 16546 24861
rect 20366 24861 20367 25039
rect 20545 24861 20546 25039
rect 24366 25039 24546 25040
rect 23734 24984 23740 24990
rect 23780 24984 23786 24990
rect 23728 24978 23734 24984
rect 23786 24978 23792 24984
rect 23728 24928 23734 24934
rect 23786 24928 23792 24934
rect 23734 24922 23740 24928
rect 23780 24922 23786 24928
rect 20366 24860 20546 24861
rect 24366 24861 24367 25039
rect 24545 24861 24546 25039
rect 28366 25039 28546 25040
rect 27734 24984 27740 24990
rect 27780 24984 27786 24990
rect 27728 24978 27734 24984
rect 27786 24978 27792 24984
rect 27728 24928 27734 24934
rect 27786 24928 27792 24934
rect 27734 24922 27740 24928
rect 27780 24922 27786 24928
rect 24366 24860 24546 24861
rect 28366 24861 28367 25039
rect 28545 24861 28546 25039
rect 32366 25039 32546 25040
rect 31734 24984 31740 24990
rect 31780 24984 31786 24990
rect 31728 24978 31734 24984
rect 31786 24978 31792 24984
rect 31728 24928 31734 24934
rect 31786 24928 31792 24934
rect 31734 24922 31740 24928
rect 31780 24922 31786 24928
rect 28366 24860 28546 24861
rect 32366 24861 32367 25039
rect 32545 24861 32546 25039
rect 36366 25039 36546 25040
rect 35734 24984 35740 24990
rect 35780 24984 35786 24990
rect 35728 24978 35734 24984
rect 35786 24978 35792 24984
rect 35728 24928 35734 24934
rect 35786 24928 35792 24934
rect 35734 24922 35740 24928
rect 35780 24922 35786 24928
rect 32366 24860 32546 24861
rect 36366 24861 36367 25039
rect 36545 24861 36546 25039
rect 39734 24984 39740 24990
rect 39780 24984 39786 24990
rect 39728 24978 39734 24984
rect 39786 24978 39792 24984
rect 39728 24928 39734 24934
rect 39786 24928 39792 24934
rect 39734 24922 39740 24928
rect 39780 24922 39786 24928
rect 36366 24860 36546 24861
rect 3262 24808 3268 24814
rect 3308 24808 3314 24814
rect 7262 24808 7268 24814
rect 7308 24808 7314 24814
rect 11262 24808 11268 24814
rect 11308 24808 11314 24814
rect 15262 24808 15268 24814
rect 15308 24808 15314 24814
rect 19262 24808 19268 24814
rect 19308 24808 19314 24814
rect 23262 24808 23268 24814
rect 23308 24808 23314 24814
rect 27262 24808 27268 24814
rect 27308 24808 27314 24814
rect 31262 24808 31268 24814
rect 31308 24808 31314 24814
rect 35262 24808 35268 24814
rect 35308 24808 35314 24814
rect 39262 24808 39268 24814
rect 39308 24808 39314 24814
rect 3256 24802 3262 24808
rect 3314 24802 3320 24808
rect 7256 24802 7262 24808
rect 7314 24802 7320 24808
rect 11256 24802 11262 24808
rect 11314 24802 11320 24808
rect 15256 24802 15262 24808
rect 15314 24802 15320 24808
rect 19256 24802 19262 24808
rect 19314 24802 19320 24808
rect 23256 24802 23262 24808
rect 23314 24802 23320 24808
rect 27256 24802 27262 24808
rect 27314 24802 27320 24808
rect 31256 24802 31262 24808
rect 31314 24802 31320 24808
rect 35256 24802 35262 24808
rect 35314 24802 35320 24808
rect 39256 24802 39262 24808
rect 39314 24802 39320 24808
rect 3256 24756 3262 24762
rect 3314 24756 3320 24762
rect 7256 24756 7262 24762
rect 7314 24756 7320 24762
rect 11256 24756 11262 24762
rect 11314 24756 11320 24762
rect 15256 24756 15262 24762
rect 15314 24756 15320 24762
rect 19256 24756 19262 24762
rect 19314 24756 19320 24762
rect 23256 24756 23262 24762
rect 23314 24756 23320 24762
rect 27256 24756 27262 24762
rect 27314 24756 27320 24762
rect 31256 24756 31262 24762
rect 31314 24756 31320 24762
rect 35256 24756 35262 24762
rect 35314 24756 35320 24762
rect 39256 24756 39262 24762
rect 39314 24756 39320 24762
rect 3262 24750 3268 24756
rect 3308 24750 3314 24756
rect 7262 24750 7268 24756
rect 7308 24750 7314 24756
rect 11262 24750 11268 24756
rect 11308 24750 11314 24756
rect 15262 24750 15268 24756
rect 15308 24750 15314 24756
rect 19262 24750 19268 24756
rect 19308 24750 19314 24756
rect 23262 24750 23268 24756
rect 23308 24750 23314 24756
rect 27262 24750 27268 24756
rect 27308 24750 27314 24756
rect 31262 24750 31268 24756
rect 31308 24750 31314 24756
rect 35262 24750 35268 24756
rect 35308 24750 35314 24756
rect 39262 24750 39268 24756
rect 39308 24750 39314 24756
rect 2386 24296 2626 24320
rect 2386 24104 2410 24296
rect 2602 24104 2626 24296
rect 2386 24080 2626 24104
rect 6386 24296 6626 24320
rect 6386 24104 6410 24296
rect 6602 24104 6626 24296
rect 6386 24080 6626 24104
rect 10386 24296 10626 24320
rect 10386 24104 10410 24296
rect 10602 24104 10626 24296
rect 10386 24080 10626 24104
rect 14386 24296 14626 24320
rect 14386 24104 14410 24296
rect 14602 24104 14626 24296
rect 14386 24080 14626 24104
rect 18386 24296 18626 24320
rect 18386 24104 18410 24296
rect 18602 24104 18626 24296
rect 18386 24080 18626 24104
rect 22386 24296 22626 24320
rect 22386 24104 22410 24296
rect 22602 24104 22626 24296
rect 22386 24080 22626 24104
rect 26386 24296 26626 24320
rect 26386 24104 26410 24296
rect 26602 24104 26626 24296
rect 26386 24080 26626 24104
rect 30386 24296 30626 24320
rect 30386 24104 30410 24296
rect 30602 24104 30626 24296
rect 30386 24080 30626 24104
rect 34386 24296 34626 24320
rect 34386 24104 34410 24296
rect 34602 24104 34626 24296
rect 34386 24080 34626 24104
rect 38386 24296 38626 24320
rect 38386 24104 38410 24296
rect 38602 24104 38626 24296
rect 38386 24080 38626 24104
rect 1982 23160 2302 23230
rect 366 22916 606 22940
rect 366 22724 390 22916
rect 582 22724 606 22916
rect 1982 22920 2006 23160
rect 2232 22920 2246 23160
rect 2256 22920 2302 23160
rect 5982 23160 6302 23230
rect 1982 22896 2302 22920
rect 4366 22916 4606 22940
rect 366 22700 606 22724
rect 4366 22724 4390 22916
rect 4582 22724 4606 22916
rect 5982 22920 6006 23160
rect 6232 22920 6246 23160
rect 6256 22920 6302 23160
rect 9982 23160 10302 23230
rect 5982 22896 6302 22920
rect 8366 22916 8606 22940
rect 2852 22709 2996 22714
rect 2852 22639 2857 22709
rect 2991 22639 2996 22709
rect 4366 22700 4606 22724
rect 8366 22724 8390 22916
rect 8582 22724 8606 22916
rect 9982 22920 10006 23160
rect 10232 22920 10246 23160
rect 10256 22920 10302 23160
rect 13982 23160 14302 23230
rect 9982 22896 10302 22920
rect 12366 22916 12606 22940
rect 6852 22709 6996 22714
rect 2852 22634 2996 22639
rect 6852 22639 6857 22709
rect 6991 22639 6996 22709
rect 8366 22700 8606 22724
rect 12366 22724 12390 22916
rect 12582 22724 12606 22916
rect 13982 22920 14006 23160
rect 14232 22920 14246 23160
rect 14256 22920 14302 23160
rect 17982 23160 18302 23230
rect 13982 22896 14302 22920
rect 16366 22916 16606 22940
rect 10852 22709 10996 22714
rect 6852 22634 6996 22639
rect 10852 22639 10857 22709
rect 10991 22639 10996 22709
rect 12366 22700 12606 22724
rect 16366 22724 16390 22916
rect 16582 22724 16606 22916
rect 17982 22920 18006 23160
rect 18232 22920 18246 23160
rect 18256 22920 18302 23160
rect 21982 23160 22302 23230
rect 17982 22896 18302 22920
rect 20366 22916 20606 22940
rect 14852 22709 14996 22714
rect 10852 22634 10996 22639
rect 14852 22639 14857 22709
rect 14991 22639 14996 22709
rect 16366 22700 16606 22724
rect 20366 22724 20390 22916
rect 20582 22724 20606 22916
rect 21982 22920 22006 23160
rect 22232 22920 22246 23160
rect 22256 22920 22302 23160
rect 25982 23160 26302 23230
rect 21982 22896 22302 22920
rect 24366 22916 24606 22940
rect 18852 22709 18996 22714
rect 14852 22634 14996 22639
rect 18852 22639 18857 22709
rect 18991 22639 18996 22709
rect 20366 22700 20606 22724
rect 24366 22724 24390 22916
rect 24582 22724 24606 22916
rect 25982 22920 26006 23160
rect 26232 22920 26246 23160
rect 26256 22920 26302 23160
rect 29982 23160 30302 23230
rect 25982 22896 26302 22920
rect 28366 22916 28606 22940
rect 22852 22709 22996 22714
rect 18852 22634 18996 22639
rect 22852 22639 22857 22709
rect 22991 22639 22996 22709
rect 24366 22700 24606 22724
rect 28366 22724 28390 22916
rect 28582 22724 28606 22916
rect 29982 22920 30006 23160
rect 30232 22920 30246 23160
rect 30256 22920 30302 23160
rect 33982 23160 34302 23230
rect 29982 22896 30302 22920
rect 32366 22916 32606 22940
rect 26852 22709 26996 22714
rect 22852 22634 22996 22639
rect 26852 22639 26857 22709
rect 26991 22639 26996 22709
rect 28366 22700 28606 22724
rect 32366 22724 32390 22916
rect 32582 22724 32606 22916
rect 33982 22920 34006 23160
rect 34232 22920 34246 23160
rect 34256 22920 34302 23160
rect 37982 23160 38302 23230
rect 33982 22896 34302 22920
rect 36366 22916 36606 22940
rect 30852 22709 30996 22714
rect 26852 22634 26996 22639
rect 30852 22639 30857 22709
rect 30991 22639 30996 22709
rect 32366 22700 32606 22724
rect 36366 22724 36390 22916
rect 36582 22724 36606 22916
rect 37982 22920 38006 23160
rect 38232 22920 38246 23160
rect 38256 22920 38302 23160
rect 37982 22896 38302 22920
rect 34852 22709 34996 22714
rect 30852 22634 30996 22639
rect 34852 22639 34857 22709
rect 34991 22639 34996 22709
rect 36366 22700 36606 22724
rect 38852 22709 38996 22714
rect 34852 22634 34996 22639
rect 38852 22639 38857 22709
rect 38991 22639 38996 22709
rect 38852 22634 38996 22639
rect 2366 22559 2546 22560
rect 2366 22381 2367 22559
rect 2545 22381 2546 22559
rect 2366 22380 2546 22381
rect 6366 22559 6546 22560
rect 6366 22381 6367 22559
rect 6545 22381 6546 22559
rect 6366 22380 6546 22381
rect 10366 22559 10546 22560
rect 10366 22381 10367 22559
rect 10545 22381 10546 22559
rect 10366 22380 10546 22381
rect 14366 22559 14546 22560
rect 14366 22381 14367 22559
rect 14545 22381 14546 22559
rect 14366 22380 14546 22381
rect 18366 22559 18546 22560
rect 18366 22381 18367 22559
rect 18545 22381 18546 22559
rect 18366 22380 18546 22381
rect 22366 22559 22546 22560
rect 22366 22381 22367 22559
rect 22545 22381 22546 22559
rect 22366 22380 22546 22381
rect 26366 22559 26546 22560
rect 26366 22381 26367 22559
rect 26545 22381 26546 22559
rect 26366 22380 26546 22381
rect 30366 22559 30546 22560
rect 30366 22381 30367 22559
rect 30545 22381 30546 22559
rect 30366 22380 30546 22381
rect 34366 22559 34546 22560
rect 34366 22381 34367 22559
rect 34545 22381 34546 22559
rect 34366 22380 34546 22381
rect 38366 22559 38546 22560
rect 38366 22381 38367 22559
rect 38545 22381 38546 22559
rect 38366 22380 38546 22381
rect 366 22039 546 22040
rect 366 21861 367 22039
rect 545 21861 546 22039
rect 4366 22039 4546 22040
rect 3734 21984 3740 21990
rect 3780 21984 3786 21990
rect 3728 21978 3734 21984
rect 3786 21978 3792 21984
rect 3728 21928 3734 21934
rect 3786 21928 3792 21934
rect 3734 21922 3740 21928
rect 3780 21922 3786 21928
rect 366 21860 546 21861
rect 4366 21861 4367 22039
rect 4545 21861 4546 22039
rect 8366 22039 8546 22040
rect 7734 21984 7740 21990
rect 7780 21984 7786 21990
rect 7728 21978 7734 21984
rect 7786 21978 7792 21984
rect 7728 21928 7734 21934
rect 7786 21928 7792 21934
rect 7734 21922 7740 21928
rect 7780 21922 7786 21928
rect 4366 21860 4546 21861
rect 8366 21861 8367 22039
rect 8545 21861 8546 22039
rect 12366 22039 12546 22040
rect 11734 21984 11740 21990
rect 11780 21984 11786 21990
rect 11728 21978 11734 21984
rect 11786 21978 11792 21984
rect 11728 21928 11734 21934
rect 11786 21928 11792 21934
rect 11734 21922 11740 21928
rect 11780 21922 11786 21928
rect 8366 21860 8546 21861
rect 12366 21861 12367 22039
rect 12545 21861 12546 22039
rect 16366 22039 16546 22040
rect 15734 21984 15740 21990
rect 15780 21984 15786 21990
rect 15728 21978 15734 21984
rect 15786 21978 15792 21984
rect 15728 21928 15734 21934
rect 15786 21928 15792 21934
rect 15734 21922 15740 21928
rect 15780 21922 15786 21928
rect 12366 21860 12546 21861
rect 16366 21861 16367 22039
rect 16545 21861 16546 22039
rect 20366 22039 20546 22040
rect 19734 21984 19740 21990
rect 19780 21984 19786 21990
rect 19728 21978 19734 21984
rect 19786 21978 19792 21984
rect 19728 21928 19734 21934
rect 19786 21928 19792 21934
rect 19734 21922 19740 21928
rect 19780 21922 19786 21928
rect 16366 21860 16546 21861
rect 20366 21861 20367 22039
rect 20545 21861 20546 22039
rect 24366 22039 24546 22040
rect 23734 21984 23740 21990
rect 23780 21984 23786 21990
rect 23728 21978 23734 21984
rect 23786 21978 23792 21984
rect 23728 21928 23734 21934
rect 23786 21928 23792 21934
rect 23734 21922 23740 21928
rect 23780 21922 23786 21928
rect 20366 21860 20546 21861
rect 24366 21861 24367 22039
rect 24545 21861 24546 22039
rect 28366 22039 28546 22040
rect 27734 21984 27740 21990
rect 27780 21984 27786 21990
rect 27728 21978 27734 21984
rect 27786 21978 27792 21984
rect 27728 21928 27734 21934
rect 27786 21928 27792 21934
rect 27734 21922 27740 21928
rect 27780 21922 27786 21928
rect 24366 21860 24546 21861
rect 28366 21861 28367 22039
rect 28545 21861 28546 22039
rect 32366 22039 32546 22040
rect 31734 21984 31740 21990
rect 31780 21984 31786 21990
rect 31728 21978 31734 21984
rect 31786 21978 31792 21984
rect 31728 21928 31734 21934
rect 31786 21928 31792 21934
rect 31734 21922 31740 21928
rect 31780 21922 31786 21928
rect 28366 21860 28546 21861
rect 32366 21861 32367 22039
rect 32545 21861 32546 22039
rect 36366 22039 36546 22040
rect 35734 21984 35740 21990
rect 35780 21984 35786 21990
rect 35728 21978 35734 21984
rect 35786 21978 35792 21984
rect 35728 21928 35734 21934
rect 35786 21928 35792 21934
rect 35734 21922 35740 21928
rect 35780 21922 35786 21928
rect 32366 21860 32546 21861
rect 36366 21861 36367 22039
rect 36545 21861 36546 22039
rect 39734 21984 39740 21990
rect 39780 21984 39786 21990
rect 39728 21978 39734 21984
rect 39786 21978 39792 21984
rect 39728 21928 39734 21934
rect 39786 21928 39792 21934
rect 39734 21922 39740 21928
rect 39780 21922 39786 21928
rect 36366 21860 36546 21861
rect 3262 21808 3268 21814
rect 3308 21808 3314 21814
rect 7262 21808 7268 21814
rect 7308 21808 7314 21814
rect 11262 21808 11268 21814
rect 11308 21808 11314 21814
rect 15262 21808 15268 21814
rect 15308 21808 15314 21814
rect 19262 21808 19268 21814
rect 19308 21808 19314 21814
rect 23262 21808 23268 21814
rect 23308 21808 23314 21814
rect 27262 21808 27268 21814
rect 27308 21808 27314 21814
rect 31262 21808 31268 21814
rect 31308 21808 31314 21814
rect 35262 21808 35268 21814
rect 35308 21808 35314 21814
rect 39262 21808 39268 21814
rect 39308 21808 39314 21814
rect 3256 21802 3262 21808
rect 3314 21802 3320 21808
rect 7256 21802 7262 21808
rect 7314 21802 7320 21808
rect 11256 21802 11262 21808
rect 11314 21802 11320 21808
rect 15256 21802 15262 21808
rect 15314 21802 15320 21808
rect 19256 21802 19262 21808
rect 19314 21802 19320 21808
rect 23256 21802 23262 21808
rect 23314 21802 23320 21808
rect 27256 21802 27262 21808
rect 27314 21802 27320 21808
rect 31256 21802 31262 21808
rect 31314 21802 31320 21808
rect 35256 21802 35262 21808
rect 35314 21802 35320 21808
rect 39256 21802 39262 21808
rect 39314 21802 39320 21808
rect 3256 21756 3262 21762
rect 3314 21756 3320 21762
rect 7256 21756 7262 21762
rect 7314 21756 7320 21762
rect 11256 21756 11262 21762
rect 11314 21756 11320 21762
rect 15256 21756 15262 21762
rect 15314 21756 15320 21762
rect 19256 21756 19262 21762
rect 19314 21756 19320 21762
rect 23256 21756 23262 21762
rect 23314 21756 23320 21762
rect 27256 21756 27262 21762
rect 27314 21756 27320 21762
rect 31256 21756 31262 21762
rect 31314 21756 31320 21762
rect 35256 21756 35262 21762
rect 35314 21756 35320 21762
rect 39256 21756 39262 21762
rect 39314 21756 39320 21762
rect 3262 21750 3268 21756
rect 3308 21750 3314 21756
rect 7262 21750 7268 21756
rect 7308 21750 7314 21756
rect 11262 21750 11268 21756
rect 11308 21750 11314 21756
rect 15262 21750 15268 21756
rect 15308 21750 15314 21756
rect 19262 21750 19268 21756
rect 19308 21750 19314 21756
rect 23262 21750 23268 21756
rect 23308 21750 23314 21756
rect 27262 21750 27268 21756
rect 27308 21750 27314 21756
rect 31262 21750 31268 21756
rect 31308 21750 31314 21756
rect 35262 21750 35268 21756
rect 35308 21750 35314 21756
rect 39262 21750 39268 21756
rect 39308 21750 39314 21756
rect 2386 21296 2626 21320
rect 2386 21104 2410 21296
rect 2602 21104 2626 21296
rect 2386 21080 2626 21104
rect 6386 21296 6626 21320
rect 6386 21104 6410 21296
rect 6602 21104 6626 21296
rect 6386 21080 6626 21104
rect 10386 21296 10626 21320
rect 10386 21104 10410 21296
rect 10602 21104 10626 21296
rect 10386 21080 10626 21104
rect 14386 21296 14626 21320
rect 14386 21104 14410 21296
rect 14602 21104 14626 21296
rect 14386 21080 14626 21104
rect 18386 21296 18626 21320
rect 18386 21104 18410 21296
rect 18602 21104 18626 21296
rect 18386 21080 18626 21104
rect 22386 21296 22626 21320
rect 22386 21104 22410 21296
rect 22602 21104 22626 21296
rect 22386 21080 22626 21104
rect 26386 21296 26626 21320
rect 26386 21104 26410 21296
rect 26602 21104 26626 21296
rect 26386 21080 26626 21104
rect 30386 21296 30626 21320
rect 30386 21104 30410 21296
rect 30602 21104 30626 21296
rect 30386 21080 30626 21104
rect 34386 21296 34626 21320
rect 34386 21104 34410 21296
rect 34602 21104 34626 21296
rect 34386 21080 34626 21104
rect 38386 21296 38626 21320
rect 38386 21104 38410 21296
rect 38602 21104 38626 21296
rect 38386 21080 38626 21104
rect 1982 20160 2302 20230
rect 366 19916 606 19940
rect 366 19724 390 19916
rect 582 19724 606 19916
rect 1982 19920 2006 20160
rect 2232 19920 2246 20160
rect 2256 19920 2302 20160
rect 5982 20160 6302 20230
rect 1982 19896 2302 19920
rect 4366 19916 4606 19940
rect 366 19700 606 19724
rect 4366 19724 4390 19916
rect 4582 19724 4606 19916
rect 5982 19920 6006 20160
rect 6232 19920 6246 20160
rect 6256 19920 6302 20160
rect 9982 20160 10302 20230
rect 5982 19896 6302 19920
rect 8366 19916 8606 19940
rect 2852 19709 2996 19714
rect 2852 19639 2857 19709
rect 2991 19639 2996 19709
rect 4366 19700 4606 19724
rect 8366 19724 8390 19916
rect 8582 19724 8606 19916
rect 9982 19920 10006 20160
rect 10232 19920 10246 20160
rect 10256 19920 10302 20160
rect 13982 20160 14302 20230
rect 9982 19896 10302 19920
rect 12366 19916 12606 19940
rect 6852 19709 6996 19714
rect 2852 19634 2996 19639
rect 6852 19639 6857 19709
rect 6991 19639 6996 19709
rect 8366 19700 8606 19724
rect 12366 19724 12390 19916
rect 12582 19724 12606 19916
rect 13982 19920 14006 20160
rect 14232 19920 14246 20160
rect 14256 19920 14302 20160
rect 17982 20160 18302 20230
rect 13982 19896 14302 19920
rect 16366 19916 16606 19940
rect 10852 19709 10996 19714
rect 6852 19634 6996 19639
rect 10852 19639 10857 19709
rect 10991 19639 10996 19709
rect 12366 19700 12606 19724
rect 16366 19724 16390 19916
rect 16582 19724 16606 19916
rect 17982 19920 18006 20160
rect 18232 19920 18246 20160
rect 18256 19920 18302 20160
rect 21982 20160 22302 20230
rect 17982 19896 18302 19920
rect 20366 19916 20606 19940
rect 14852 19709 14996 19714
rect 10852 19634 10996 19639
rect 14852 19639 14857 19709
rect 14991 19639 14996 19709
rect 16366 19700 16606 19724
rect 20366 19724 20390 19916
rect 20582 19724 20606 19916
rect 21982 19920 22006 20160
rect 22232 19920 22246 20160
rect 22256 19920 22302 20160
rect 25982 20160 26302 20230
rect 21982 19896 22302 19920
rect 24366 19916 24606 19940
rect 18852 19709 18996 19714
rect 14852 19634 14996 19639
rect 18852 19639 18857 19709
rect 18991 19639 18996 19709
rect 20366 19700 20606 19724
rect 24366 19724 24390 19916
rect 24582 19724 24606 19916
rect 25982 19920 26006 20160
rect 26232 19920 26246 20160
rect 26256 19920 26302 20160
rect 29982 20160 30302 20230
rect 25982 19896 26302 19920
rect 28366 19916 28606 19940
rect 22852 19709 22996 19714
rect 18852 19634 18996 19639
rect 22852 19639 22857 19709
rect 22991 19639 22996 19709
rect 24366 19700 24606 19724
rect 28366 19724 28390 19916
rect 28582 19724 28606 19916
rect 29982 19920 30006 20160
rect 30232 19920 30246 20160
rect 30256 19920 30302 20160
rect 33982 20160 34302 20230
rect 29982 19896 30302 19920
rect 32366 19916 32606 19940
rect 26852 19709 26996 19714
rect 22852 19634 22996 19639
rect 26852 19639 26857 19709
rect 26991 19639 26996 19709
rect 28366 19700 28606 19724
rect 32366 19724 32390 19916
rect 32582 19724 32606 19916
rect 33982 19920 34006 20160
rect 34232 19920 34246 20160
rect 34256 19920 34302 20160
rect 37982 20160 38302 20230
rect 33982 19896 34302 19920
rect 36366 19916 36606 19940
rect 30852 19709 30996 19714
rect 26852 19634 26996 19639
rect 30852 19639 30857 19709
rect 30991 19639 30996 19709
rect 32366 19700 32606 19724
rect 36366 19724 36390 19916
rect 36582 19724 36606 19916
rect 37982 19920 38006 20160
rect 38232 19920 38246 20160
rect 38256 19920 38302 20160
rect 37982 19896 38302 19920
rect 34852 19709 34996 19714
rect 30852 19634 30996 19639
rect 34852 19639 34857 19709
rect 34991 19639 34996 19709
rect 36366 19700 36606 19724
rect 38852 19709 38996 19714
rect 34852 19634 34996 19639
rect 38852 19639 38857 19709
rect 38991 19639 38996 19709
rect 38852 19634 38996 19639
rect 2366 19559 2546 19560
rect 2366 19381 2367 19559
rect 2545 19381 2546 19559
rect 2366 19380 2546 19381
rect 6366 19559 6546 19560
rect 6366 19381 6367 19559
rect 6545 19381 6546 19559
rect 6366 19380 6546 19381
rect 10366 19559 10546 19560
rect 10366 19381 10367 19559
rect 10545 19381 10546 19559
rect 10366 19380 10546 19381
rect 14366 19559 14546 19560
rect 14366 19381 14367 19559
rect 14545 19381 14546 19559
rect 14366 19380 14546 19381
rect 18366 19559 18546 19560
rect 18366 19381 18367 19559
rect 18545 19381 18546 19559
rect 18366 19380 18546 19381
rect 22366 19559 22546 19560
rect 22366 19381 22367 19559
rect 22545 19381 22546 19559
rect 22366 19380 22546 19381
rect 26366 19559 26546 19560
rect 26366 19381 26367 19559
rect 26545 19381 26546 19559
rect 26366 19380 26546 19381
rect 30366 19559 30546 19560
rect 30366 19381 30367 19559
rect 30545 19381 30546 19559
rect 30366 19380 30546 19381
rect 34366 19559 34546 19560
rect 34366 19381 34367 19559
rect 34545 19381 34546 19559
rect 34366 19380 34546 19381
rect 38366 19559 38546 19560
rect 38366 19381 38367 19559
rect 38545 19381 38546 19559
rect 38366 19380 38546 19381
rect 366 19039 546 19040
rect 366 18861 367 19039
rect 545 18861 546 19039
rect 4366 19039 4546 19040
rect 3734 18984 3740 18990
rect 3780 18984 3786 18990
rect 3728 18978 3734 18984
rect 3786 18978 3792 18984
rect 3728 18928 3734 18934
rect 3786 18928 3792 18934
rect 3734 18922 3740 18928
rect 3780 18922 3786 18928
rect 366 18860 546 18861
rect 4366 18861 4367 19039
rect 4545 18861 4546 19039
rect 8366 19039 8546 19040
rect 7734 18984 7740 18990
rect 7780 18984 7786 18990
rect 7728 18978 7734 18984
rect 7786 18978 7792 18984
rect 7728 18928 7734 18934
rect 7786 18928 7792 18934
rect 7734 18922 7740 18928
rect 7780 18922 7786 18928
rect 4366 18860 4546 18861
rect 8366 18861 8367 19039
rect 8545 18861 8546 19039
rect 12366 19039 12546 19040
rect 11734 18984 11740 18990
rect 11780 18984 11786 18990
rect 11728 18978 11734 18984
rect 11786 18978 11792 18984
rect 11728 18928 11734 18934
rect 11786 18928 11792 18934
rect 11734 18922 11740 18928
rect 11780 18922 11786 18928
rect 8366 18860 8546 18861
rect 12366 18861 12367 19039
rect 12545 18861 12546 19039
rect 16366 19039 16546 19040
rect 15734 18984 15740 18990
rect 15780 18984 15786 18990
rect 15728 18978 15734 18984
rect 15786 18978 15792 18984
rect 15728 18928 15734 18934
rect 15786 18928 15792 18934
rect 15734 18922 15740 18928
rect 15780 18922 15786 18928
rect 12366 18860 12546 18861
rect 16366 18861 16367 19039
rect 16545 18861 16546 19039
rect 20366 19039 20546 19040
rect 19734 18984 19740 18990
rect 19780 18984 19786 18990
rect 19728 18978 19734 18984
rect 19786 18978 19792 18984
rect 19728 18928 19734 18934
rect 19786 18928 19792 18934
rect 19734 18922 19740 18928
rect 19780 18922 19786 18928
rect 16366 18860 16546 18861
rect 20366 18861 20367 19039
rect 20545 18861 20546 19039
rect 24366 19039 24546 19040
rect 23734 18984 23740 18990
rect 23780 18984 23786 18990
rect 23728 18978 23734 18984
rect 23786 18978 23792 18984
rect 23728 18928 23734 18934
rect 23786 18928 23792 18934
rect 23734 18922 23740 18928
rect 23780 18922 23786 18928
rect 20366 18860 20546 18861
rect 24366 18861 24367 19039
rect 24545 18861 24546 19039
rect 28366 19039 28546 19040
rect 27734 18984 27740 18990
rect 27780 18984 27786 18990
rect 27728 18978 27734 18984
rect 27786 18978 27792 18984
rect 27728 18928 27734 18934
rect 27786 18928 27792 18934
rect 27734 18922 27740 18928
rect 27780 18922 27786 18928
rect 24366 18860 24546 18861
rect 28366 18861 28367 19039
rect 28545 18861 28546 19039
rect 32366 19039 32546 19040
rect 31734 18984 31740 18990
rect 31780 18984 31786 18990
rect 31728 18978 31734 18984
rect 31786 18978 31792 18984
rect 31728 18928 31734 18934
rect 31786 18928 31792 18934
rect 31734 18922 31740 18928
rect 31780 18922 31786 18928
rect 28366 18860 28546 18861
rect 32366 18861 32367 19039
rect 32545 18861 32546 19039
rect 36366 19039 36546 19040
rect 35734 18984 35740 18990
rect 35780 18984 35786 18990
rect 35728 18978 35734 18984
rect 35786 18978 35792 18984
rect 35728 18928 35734 18934
rect 35786 18928 35792 18934
rect 35734 18922 35740 18928
rect 35780 18922 35786 18928
rect 32366 18860 32546 18861
rect 36366 18861 36367 19039
rect 36545 18861 36546 19039
rect 39734 18984 39740 18990
rect 39780 18984 39786 18990
rect 39728 18978 39734 18984
rect 39786 18978 39792 18984
rect 39728 18928 39734 18934
rect 39786 18928 39792 18934
rect 39734 18922 39740 18928
rect 39780 18922 39786 18928
rect 36366 18860 36546 18861
rect 3262 18808 3268 18814
rect 3308 18808 3314 18814
rect 7262 18808 7268 18814
rect 7308 18808 7314 18814
rect 11262 18808 11268 18814
rect 11308 18808 11314 18814
rect 15262 18808 15268 18814
rect 15308 18808 15314 18814
rect 19262 18808 19268 18814
rect 19308 18808 19314 18814
rect 23262 18808 23268 18814
rect 23308 18808 23314 18814
rect 27262 18808 27268 18814
rect 27308 18808 27314 18814
rect 31262 18808 31268 18814
rect 31308 18808 31314 18814
rect 35262 18808 35268 18814
rect 35308 18808 35314 18814
rect 39262 18808 39268 18814
rect 39308 18808 39314 18814
rect 3256 18802 3262 18808
rect 3314 18802 3320 18808
rect 7256 18802 7262 18808
rect 7314 18802 7320 18808
rect 11256 18802 11262 18808
rect 11314 18802 11320 18808
rect 15256 18802 15262 18808
rect 15314 18802 15320 18808
rect 19256 18802 19262 18808
rect 19314 18802 19320 18808
rect 23256 18802 23262 18808
rect 23314 18802 23320 18808
rect 27256 18802 27262 18808
rect 27314 18802 27320 18808
rect 31256 18802 31262 18808
rect 31314 18802 31320 18808
rect 35256 18802 35262 18808
rect 35314 18802 35320 18808
rect 39256 18802 39262 18808
rect 39314 18802 39320 18808
rect 3256 18756 3262 18762
rect 3314 18756 3320 18762
rect 7256 18756 7262 18762
rect 7314 18756 7320 18762
rect 11256 18756 11262 18762
rect 11314 18756 11320 18762
rect 15256 18756 15262 18762
rect 15314 18756 15320 18762
rect 19256 18756 19262 18762
rect 19314 18756 19320 18762
rect 23256 18756 23262 18762
rect 23314 18756 23320 18762
rect 27256 18756 27262 18762
rect 27314 18756 27320 18762
rect 31256 18756 31262 18762
rect 31314 18756 31320 18762
rect 35256 18756 35262 18762
rect 35314 18756 35320 18762
rect 39256 18756 39262 18762
rect 39314 18756 39320 18762
rect 3262 18750 3268 18756
rect 3308 18750 3314 18756
rect 7262 18750 7268 18756
rect 7308 18750 7314 18756
rect 11262 18750 11268 18756
rect 11308 18750 11314 18756
rect 15262 18750 15268 18756
rect 15308 18750 15314 18756
rect 19262 18750 19268 18756
rect 19308 18750 19314 18756
rect 23262 18750 23268 18756
rect 23308 18750 23314 18756
rect 27262 18750 27268 18756
rect 27308 18750 27314 18756
rect 31262 18750 31268 18756
rect 31308 18750 31314 18756
rect 35262 18750 35268 18756
rect 35308 18750 35314 18756
rect 39262 18750 39268 18756
rect 39308 18750 39314 18756
rect 2386 18296 2626 18320
rect 2386 18104 2410 18296
rect 2602 18104 2626 18296
rect 2386 18080 2626 18104
rect 6386 18296 6626 18320
rect 6386 18104 6410 18296
rect 6602 18104 6626 18296
rect 6386 18080 6626 18104
rect 10386 18296 10626 18320
rect 10386 18104 10410 18296
rect 10602 18104 10626 18296
rect 10386 18080 10626 18104
rect 14386 18296 14626 18320
rect 14386 18104 14410 18296
rect 14602 18104 14626 18296
rect 14386 18080 14626 18104
rect 18386 18296 18626 18320
rect 18386 18104 18410 18296
rect 18602 18104 18626 18296
rect 18386 18080 18626 18104
rect 22386 18296 22626 18320
rect 22386 18104 22410 18296
rect 22602 18104 22626 18296
rect 22386 18080 22626 18104
rect 26386 18296 26626 18320
rect 26386 18104 26410 18296
rect 26602 18104 26626 18296
rect 26386 18080 26626 18104
rect 30386 18296 30626 18320
rect 30386 18104 30410 18296
rect 30602 18104 30626 18296
rect 30386 18080 30626 18104
rect 34386 18296 34626 18320
rect 34386 18104 34410 18296
rect 34602 18104 34626 18296
rect 34386 18080 34626 18104
rect 38386 18296 38626 18320
rect 38386 18104 38410 18296
rect 38602 18104 38626 18296
rect 38386 18080 38626 18104
rect 1982 17160 2302 17230
rect 366 16916 606 16940
rect 366 16724 390 16916
rect 582 16724 606 16916
rect 1982 16920 2006 17160
rect 2232 16920 2246 17160
rect 2256 16920 2302 17160
rect 5982 17160 6302 17230
rect 1982 16896 2302 16920
rect 4366 16916 4606 16940
rect 366 16700 606 16724
rect 4366 16724 4390 16916
rect 4582 16724 4606 16916
rect 5982 16920 6006 17160
rect 6232 16920 6246 17160
rect 6256 16920 6302 17160
rect 9982 17160 10302 17230
rect 5982 16896 6302 16920
rect 8366 16916 8606 16940
rect 2852 16709 2996 16714
rect 2852 16639 2857 16709
rect 2991 16639 2996 16709
rect 4366 16700 4606 16724
rect 8366 16724 8390 16916
rect 8582 16724 8606 16916
rect 9982 16920 10006 17160
rect 10232 16920 10246 17160
rect 10256 16920 10302 17160
rect 13982 17160 14302 17230
rect 9982 16896 10302 16920
rect 12366 16916 12606 16940
rect 6852 16709 6996 16714
rect 2852 16634 2996 16639
rect 6852 16639 6857 16709
rect 6991 16639 6996 16709
rect 8366 16700 8606 16724
rect 12366 16724 12390 16916
rect 12582 16724 12606 16916
rect 13982 16920 14006 17160
rect 14232 16920 14246 17160
rect 14256 16920 14302 17160
rect 17982 17160 18302 17230
rect 13982 16896 14302 16920
rect 16366 16916 16606 16940
rect 10852 16709 10996 16714
rect 6852 16634 6996 16639
rect 10852 16639 10857 16709
rect 10991 16639 10996 16709
rect 12366 16700 12606 16724
rect 16366 16724 16390 16916
rect 16582 16724 16606 16916
rect 17982 16920 18006 17160
rect 18232 16920 18246 17160
rect 18256 16920 18302 17160
rect 21982 17160 22302 17230
rect 17982 16896 18302 16920
rect 20366 16916 20606 16940
rect 14852 16709 14996 16714
rect 10852 16634 10996 16639
rect 14852 16639 14857 16709
rect 14991 16639 14996 16709
rect 16366 16700 16606 16724
rect 20366 16724 20390 16916
rect 20582 16724 20606 16916
rect 21982 16920 22006 17160
rect 22232 16920 22246 17160
rect 22256 16920 22302 17160
rect 25982 17160 26302 17230
rect 21982 16896 22302 16920
rect 24366 16916 24606 16940
rect 18852 16709 18996 16714
rect 14852 16634 14996 16639
rect 18852 16639 18857 16709
rect 18991 16639 18996 16709
rect 20366 16700 20606 16724
rect 24366 16724 24390 16916
rect 24582 16724 24606 16916
rect 25982 16920 26006 17160
rect 26232 16920 26246 17160
rect 26256 16920 26302 17160
rect 29982 17160 30302 17230
rect 25982 16896 26302 16920
rect 28366 16916 28606 16940
rect 22852 16709 22996 16714
rect 18852 16634 18996 16639
rect 22852 16639 22857 16709
rect 22991 16639 22996 16709
rect 24366 16700 24606 16724
rect 28366 16724 28390 16916
rect 28582 16724 28606 16916
rect 29982 16920 30006 17160
rect 30232 16920 30246 17160
rect 30256 16920 30302 17160
rect 33982 17160 34302 17230
rect 29982 16896 30302 16920
rect 32366 16916 32606 16940
rect 26852 16709 26996 16714
rect 22852 16634 22996 16639
rect 26852 16639 26857 16709
rect 26991 16639 26996 16709
rect 28366 16700 28606 16724
rect 32366 16724 32390 16916
rect 32582 16724 32606 16916
rect 33982 16920 34006 17160
rect 34232 16920 34246 17160
rect 34256 16920 34302 17160
rect 37982 17160 38302 17230
rect 33982 16896 34302 16920
rect 36366 16916 36606 16940
rect 30852 16709 30996 16714
rect 26852 16634 26996 16639
rect 30852 16639 30857 16709
rect 30991 16639 30996 16709
rect 32366 16700 32606 16724
rect 36366 16724 36390 16916
rect 36582 16724 36606 16916
rect 37982 16920 38006 17160
rect 38232 16920 38246 17160
rect 38256 16920 38302 17160
rect 37982 16896 38302 16920
rect 34852 16709 34996 16714
rect 30852 16634 30996 16639
rect 34852 16639 34857 16709
rect 34991 16639 34996 16709
rect 36366 16700 36606 16724
rect 38852 16709 38996 16714
rect 34852 16634 34996 16639
rect 38852 16639 38857 16709
rect 38991 16639 38996 16709
rect 38852 16634 38996 16639
rect 2366 16559 2546 16560
rect 2366 16381 2367 16559
rect 2545 16381 2546 16559
rect 2366 16380 2546 16381
rect 6366 16559 6546 16560
rect 6366 16381 6367 16559
rect 6545 16381 6546 16559
rect 6366 16380 6546 16381
rect 10366 16559 10546 16560
rect 10366 16381 10367 16559
rect 10545 16381 10546 16559
rect 10366 16380 10546 16381
rect 14366 16559 14546 16560
rect 14366 16381 14367 16559
rect 14545 16381 14546 16559
rect 14366 16380 14546 16381
rect 18366 16559 18546 16560
rect 18366 16381 18367 16559
rect 18545 16381 18546 16559
rect 18366 16380 18546 16381
rect 22366 16559 22546 16560
rect 22366 16381 22367 16559
rect 22545 16381 22546 16559
rect 22366 16380 22546 16381
rect 26366 16559 26546 16560
rect 26366 16381 26367 16559
rect 26545 16381 26546 16559
rect 26366 16380 26546 16381
rect 30366 16559 30546 16560
rect 30366 16381 30367 16559
rect 30545 16381 30546 16559
rect 30366 16380 30546 16381
rect 34366 16559 34546 16560
rect 34366 16381 34367 16559
rect 34545 16381 34546 16559
rect 34366 16380 34546 16381
rect 38366 16559 38546 16560
rect 38366 16381 38367 16559
rect 38545 16381 38546 16559
rect 38366 16380 38546 16381
rect 366 16039 546 16040
rect 366 15861 367 16039
rect 545 15861 546 16039
rect 4366 16039 4546 16040
rect 3734 15984 3740 15990
rect 3780 15984 3786 15990
rect 3728 15978 3734 15984
rect 3786 15978 3792 15984
rect 3728 15928 3734 15934
rect 3786 15928 3792 15934
rect 3734 15922 3740 15928
rect 3780 15922 3786 15928
rect 366 15860 546 15861
rect 4366 15861 4367 16039
rect 4545 15861 4546 16039
rect 8366 16039 8546 16040
rect 7734 15984 7740 15990
rect 7780 15984 7786 15990
rect 7728 15978 7734 15984
rect 7786 15978 7792 15984
rect 7728 15928 7734 15934
rect 7786 15928 7792 15934
rect 7734 15922 7740 15928
rect 7780 15922 7786 15928
rect 4366 15860 4546 15861
rect 8366 15861 8367 16039
rect 8545 15861 8546 16039
rect 12366 16039 12546 16040
rect 11734 15984 11740 15990
rect 11780 15984 11786 15990
rect 11728 15978 11734 15984
rect 11786 15978 11792 15984
rect 11728 15928 11734 15934
rect 11786 15928 11792 15934
rect 11734 15922 11740 15928
rect 11780 15922 11786 15928
rect 8366 15860 8546 15861
rect 12366 15861 12367 16039
rect 12545 15861 12546 16039
rect 16366 16039 16546 16040
rect 15734 15984 15740 15990
rect 15780 15984 15786 15990
rect 15728 15978 15734 15984
rect 15786 15978 15792 15984
rect 15728 15928 15734 15934
rect 15786 15928 15792 15934
rect 15734 15922 15740 15928
rect 15780 15922 15786 15928
rect 12366 15860 12546 15861
rect 16366 15861 16367 16039
rect 16545 15861 16546 16039
rect 20366 16039 20546 16040
rect 19734 15984 19740 15990
rect 19780 15984 19786 15990
rect 19728 15978 19734 15984
rect 19786 15978 19792 15984
rect 19728 15928 19734 15934
rect 19786 15928 19792 15934
rect 19734 15922 19740 15928
rect 19780 15922 19786 15928
rect 16366 15860 16546 15861
rect 20366 15861 20367 16039
rect 20545 15861 20546 16039
rect 24366 16039 24546 16040
rect 23734 15984 23740 15990
rect 23780 15984 23786 15990
rect 23728 15978 23734 15984
rect 23786 15978 23792 15984
rect 23728 15928 23734 15934
rect 23786 15928 23792 15934
rect 23734 15922 23740 15928
rect 23780 15922 23786 15928
rect 20366 15860 20546 15861
rect 24366 15861 24367 16039
rect 24545 15861 24546 16039
rect 28366 16039 28546 16040
rect 27734 15984 27740 15990
rect 27780 15984 27786 15990
rect 27728 15978 27734 15984
rect 27786 15978 27792 15984
rect 27728 15928 27734 15934
rect 27786 15928 27792 15934
rect 27734 15922 27740 15928
rect 27780 15922 27786 15928
rect 24366 15860 24546 15861
rect 28366 15861 28367 16039
rect 28545 15861 28546 16039
rect 32366 16039 32546 16040
rect 31734 15984 31740 15990
rect 31780 15984 31786 15990
rect 31728 15978 31734 15984
rect 31786 15978 31792 15984
rect 31728 15928 31734 15934
rect 31786 15928 31792 15934
rect 31734 15922 31740 15928
rect 31780 15922 31786 15928
rect 28366 15860 28546 15861
rect 32366 15861 32367 16039
rect 32545 15861 32546 16039
rect 36366 16039 36546 16040
rect 35734 15984 35740 15990
rect 35780 15984 35786 15990
rect 35728 15978 35734 15984
rect 35786 15978 35792 15984
rect 35728 15928 35734 15934
rect 35786 15928 35792 15934
rect 35734 15922 35740 15928
rect 35780 15922 35786 15928
rect 32366 15860 32546 15861
rect 36366 15861 36367 16039
rect 36545 15861 36546 16039
rect 39734 15984 39740 15990
rect 39780 15984 39786 15990
rect 39728 15978 39734 15984
rect 39786 15978 39792 15984
rect 39728 15928 39734 15934
rect 39786 15928 39792 15934
rect 39734 15922 39740 15928
rect 39780 15922 39786 15928
rect 36366 15860 36546 15861
rect 3262 15808 3268 15814
rect 3308 15808 3314 15814
rect 7262 15808 7268 15814
rect 7308 15808 7314 15814
rect 11262 15808 11268 15814
rect 11308 15808 11314 15814
rect 15262 15808 15268 15814
rect 15308 15808 15314 15814
rect 19262 15808 19268 15814
rect 19308 15808 19314 15814
rect 23262 15808 23268 15814
rect 23308 15808 23314 15814
rect 27262 15808 27268 15814
rect 27308 15808 27314 15814
rect 31262 15808 31268 15814
rect 31308 15808 31314 15814
rect 35262 15808 35268 15814
rect 35308 15808 35314 15814
rect 39262 15808 39268 15814
rect 39308 15808 39314 15814
rect 3256 15802 3262 15808
rect 3314 15802 3320 15808
rect 7256 15802 7262 15808
rect 7314 15802 7320 15808
rect 11256 15802 11262 15808
rect 11314 15802 11320 15808
rect 15256 15802 15262 15808
rect 15314 15802 15320 15808
rect 19256 15802 19262 15808
rect 19314 15802 19320 15808
rect 23256 15802 23262 15808
rect 23314 15802 23320 15808
rect 27256 15802 27262 15808
rect 27314 15802 27320 15808
rect 31256 15802 31262 15808
rect 31314 15802 31320 15808
rect 35256 15802 35262 15808
rect 35314 15802 35320 15808
rect 39256 15802 39262 15808
rect 39314 15802 39320 15808
rect 3256 15756 3262 15762
rect 3314 15756 3320 15762
rect 7256 15756 7262 15762
rect 7314 15756 7320 15762
rect 11256 15756 11262 15762
rect 11314 15756 11320 15762
rect 15256 15756 15262 15762
rect 15314 15756 15320 15762
rect 19256 15756 19262 15762
rect 19314 15756 19320 15762
rect 23256 15756 23262 15762
rect 23314 15756 23320 15762
rect 27256 15756 27262 15762
rect 27314 15756 27320 15762
rect 31256 15756 31262 15762
rect 31314 15756 31320 15762
rect 35256 15756 35262 15762
rect 35314 15756 35320 15762
rect 39256 15756 39262 15762
rect 39314 15756 39320 15762
rect 3262 15750 3268 15756
rect 3308 15750 3314 15756
rect 7262 15750 7268 15756
rect 7308 15750 7314 15756
rect 11262 15750 11268 15756
rect 11308 15750 11314 15756
rect 15262 15750 15268 15756
rect 15308 15750 15314 15756
rect 19262 15750 19268 15756
rect 19308 15750 19314 15756
rect 23262 15750 23268 15756
rect 23308 15750 23314 15756
rect 27262 15750 27268 15756
rect 27308 15750 27314 15756
rect 31262 15750 31268 15756
rect 31308 15750 31314 15756
rect 35262 15750 35268 15756
rect 35308 15750 35314 15756
rect 39262 15750 39268 15756
rect 39308 15750 39314 15756
rect 2386 15296 2626 15320
rect 2386 15104 2410 15296
rect 2602 15104 2626 15296
rect 2386 15080 2626 15104
rect 6386 15296 6626 15320
rect 6386 15104 6410 15296
rect 6602 15104 6626 15296
rect 6386 15080 6626 15104
rect 10386 15296 10626 15320
rect 10386 15104 10410 15296
rect 10602 15104 10626 15296
rect 10386 15080 10626 15104
rect 14386 15296 14626 15320
rect 14386 15104 14410 15296
rect 14602 15104 14626 15296
rect 14386 15080 14626 15104
rect 18386 15296 18626 15320
rect 18386 15104 18410 15296
rect 18602 15104 18626 15296
rect 18386 15080 18626 15104
rect 22386 15296 22626 15320
rect 22386 15104 22410 15296
rect 22602 15104 22626 15296
rect 22386 15080 22626 15104
rect 26386 15296 26626 15320
rect 26386 15104 26410 15296
rect 26602 15104 26626 15296
rect 26386 15080 26626 15104
rect 30386 15296 30626 15320
rect 30386 15104 30410 15296
rect 30602 15104 30626 15296
rect 30386 15080 30626 15104
rect 34386 15296 34626 15320
rect 34386 15104 34410 15296
rect 34602 15104 34626 15296
rect 34386 15080 34626 15104
rect 38386 15296 38626 15320
rect 38386 15104 38410 15296
rect 38602 15104 38626 15296
rect 38386 15080 38626 15104
rect 1982 14160 2302 14230
rect 366 13916 606 13940
rect 366 13724 390 13916
rect 582 13724 606 13916
rect 1982 13920 2006 14160
rect 2232 13920 2246 14160
rect 2256 13920 2302 14160
rect 5982 14160 6302 14230
rect 1982 13896 2302 13920
rect 4366 13916 4606 13940
rect 366 13700 606 13724
rect 4366 13724 4390 13916
rect 4582 13724 4606 13916
rect 5982 13920 6006 14160
rect 6232 13920 6246 14160
rect 6256 13920 6302 14160
rect 9982 14160 10302 14230
rect 5982 13896 6302 13920
rect 8366 13916 8606 13940
rect 2852 13709 2996 13714
rect 2852 13639 2857 13709
rect 2991 13639 2996 13709
rect 4366 13700 4606 13724
rect 8366 13724 8390 13916
rect 8582 13724 8606 13916
rect 9982 13920 10006 14160
rect 10232 13920 10246 14160
rect 10256 13920 10302 14160
rect 13982 14160 14302 14230
rect 9982 13896 10302 13920
rect 12366 13916 12606 13940
rect 6852 13709 6996 13714
rect 2852 13634 2996 13639
rect 6852 13639 6857 13709
rect 6991 13639 6996 13709
rect 8366 13700 8606 13724
rect 12366 13724 12390 13916
rect 12582 13724 12606 13916
rect 13982 13920 14006 14160
rect 14232 13920 14246 14160
rect 14256 13920 14302 14160
rect 17982 14160 18302 14230
rect 13982 13896 14302 13920
rect 16366 13916 16606 13940
rect 10852 13709 10996 13714
rect 6852 13634 6996 13639
rect 10852 13639 10857 13709
rect 10991 13639 10996 13709
rect 12366 13700 12606 13724
rect 16366 13724 16390 13916
rect 16582 13724 16606 13916
rect 17982 13920 18006 14160
rect 18232 13920 18246 14160
rect 18256 13920 18302 14160
rect 21982 14160 22302 14230
rect 17982 13896 18302 13920
rect 20366 13916 20606 13940
rect 14852 13709 14996 13714
rect 10852 13634 10996 13639
rect 14852 13639 14857 13709
rect 14991 13639 14996 13709
rect 16366 13700 16606 13724
rect 20366 13724 20390 13916
rect 20582 13724 20606 13916
rect 21982 13920 22006 14160
rect 22232 13920 22246 14160
rect 22256 13920 22302 14160
rect 25982 14160 26302 14230
rect 21982 13896 22302 13920
rect 24366 13916 24606 13940
rect 18852 13709 18996 13714
rect 14852 13634 14996 13639
rect 18852 13639 18857 13709
rect 18991 13639 18996 13709
rect 20366 13700 20606 13724
rect 24366 13724 24390 13916
rect 24582 13724 24606 13916
rect 25982 13920 26006 14160
rect 26232 13920 26246 14160
rect 26256 13920 26302 14160
rect 29982 14160 30302 14230
rect 25982 13896 26302 13920
rect 28366 13916 28606 13940
rect 22852 13709 22996 13714
rect 18852 13634 18996 13639
rect 22852 13639 22857 13709
rect 22991 13639 22996 13709
rect 24366 13700 24606 13724
rect 28366 13724 28390 13916
rect 28582 13724 28606 13916
rect 29982 13920 30006 14160
rect 30232 13920 30246 14160
rect 30256 13920 30302 14160
rect 33982 14160 34302 14230
rect 29982 13896 30302 13920
rect 32366 13916 32606 13940
rect 26852 13709 26996 13714
rect 22852 13634 22996 13639
rect 26852 13639 26857 13709
rect 26991 13639 26996 13709
rect 28366 13700 28606 13724
rect 32366 13724 32390 13916
rect 32582 13724 32606 13916
rect 33982 13920 34006 14160
rect 34232 13920 34246 14160
rect 34256 13920 34302 14160
rect 37982 14160 38302 14230
rect 33982 13896 34302 13920
rect 36366 13916 36606 13940
rect 30852 13709 30996 13714
rect 26852 13634 26996 13639
rect 30852 13639 30857 13709
rect 30991 13639 30996 13709
rect 32366 13700 32606 13724
rect 36366 13724 36390 13916
rect 36582 13724 36606 13916
rect 37982 13920 38006 14160
rect 38232 13920 38246 14160
rect 38256 13920 38302 14160
rect 37982 13896 38302 13920
rect 34852 13709 34996 13714
rect 30852 13634 30996 13639
rect 34852 13639 34857 13709
rect 34991 13639 34996 13709
rect 36366 13700 36606 13724
rect 38852 13709 38996 13714
rect 34852 13634 34996 13639
rect 38852 13639 38857 13709
rect 38991 13639 38996 13709
rect 38852 13634 38996 13639
rect 2366 13559 2546 13560
rect 2366 13381 2367 13559
rect 2545 13381 2546 13559
rect 2366 13380 2546 13381
rect 6366 13559 6546 13560
rect 6366 13381 6367 13559
rect 6545 13381 6546 13559
rect 6366 13380 6546 13381
rect 10366 13559 10546 13560
rect 10366 13381 10367 13559
rect 10545 13381 10546 13559
rect 10366 13380 10546 13381
rect 14366 13559 14546 13560
rect 14366 13381 14367 13559
rect 14545 13381 14546 13559
rect 14366 13380 14546 13381
rect 18366 13559 18546 13560
rect 18366 13381 18367 13559
rect 18545 13381 18546 13559
rect 18366 13380 18546 13381
rect 22366 13559 22546 13560
rect 22366 13381 22367 13559
rect 22545 13381 22546 13559
rect 22366 13380 22546 13381
rect 26366 13559 26546 13560
rect 26366 13381 26367 13559
rect 26545 13381 26546 13559
rect 26366 13380 26546 13381
rect 30366 13559 30546 13560
rect 30366 13381 30367 13559
rect 30545 13381 30546 13559
rect 30366 13380 30546 13381
rect 34366 13559 34546 13560
rect 34366 13381 34367 13559
rect 34545 13381 34546 13559
rect 34366 13380 34546 13381
rect 38366 13559 38546 13560
rect 38366 13381 38367 13559
rect 38545 13381 38546 13559
rect 38366 13380 38546 13381
rect 366 13039 546 13040
rect 366 12861 367 13039
rect 545 12861 546 13039
rect 4366 13039 4546 13040
rect 3734 12984 3740 12990
rect 3780 12984 3786 12990
rect 3728 12978 3734 12984
rect 3786 12978 3792 12984
rect 3728 12928 3734 12934
rect 3786 12928 3792 12934
rect 3734 12922 3740 12928
rect 3780 12922 3786 12928
rect 366 12860 546 12861
rect 4366 12861 4367 13039
rect 4545 12861 4546 13039
rect 8366 13039 8546 13040
rect 7734 12984 7740 12990
rect 7780 12984 7786 12990
rect 7728 12978 7734 12984
rect 7786 12978 7792 12984
rect 7728 12928 7734 12934
rect 7786 12928 7792 12934
rect 7734 12922 7740 12928
rect 7780 12922 7786 12928
rect 4366 12860 4546 12861
rect 8366 12861 8367 13039
rect 8545 12861 8546 13039
rect 12366 13039 12546 13040
rect 11734 12984 11740 12990
rect 11780 12984 11786 12990
rect 11728 12978 11734 12984
rect 11786 12978 11792 12984
rect 11728 12928 11734 12934
rect 11786 12928 11792 12934
rect 11734 12922 11740 12928
rect 11780 12922 11786 12928
rect 8366 12860 8546 12861
rect 12366 12861 12367 13039
rect 12545 12861 12546 13039
rect 16366 13039 16546 13040
rect 15734 12984 15740 12990
rect 15780 12984 15786 12990
rect 15728 12978 15734 12984
rect 15786 12978 15792 12984
rect 15728 12928 15734 12934
rect 15786 12928 15792 12934
rect 15734 12922 15740 12928
rect 15780 12922 15786 12928
rect 12366 12860 12546 12861
rect 16366 12861 16367 13039
rect 16545 12861 16546 13039
rect 20366 13039 20546 13040
rect 19734 12984 19740 12990
rect 19780 12984 19786 12990
rect 19728 12978 19734 12984
rect 19786 12978 19792 12984
rect 19728 12928 19734 12934
rect 19786 12928 19792 12934
rect 19734 12922 19740 12928
rect 19780 12922 19786 12928
rect 16366 12860 16546 12861
rect 20366 12861 20367 13039
rect 20545 12861 20546 13039
rect 24366 13039 24546 13040
rect 23734 12984 23740 12990
rect 23780 12984 23786 12990
rect 23728 12978 23734 12984
rect 23786 12978 23792 12984
rect 23728 12928 23734 12934
rect 23786 12928 23792 12934
rect 23734 12922 23740 12928
rect 23780 12922 23786 12928
rect 20366 12860 20546 12861
rect 24366 12861 24367 13039
rect 24545 12861 24546 13039
rect 28366 13039 28546 13040
rect 27734 12984 27740 12990
rect 27780 12984 27786 12990
rect 27728 12978 27734 12984
rect 27786 12978 27792 12984
rect 27728 12928 27734 12934
rect 27786 12928 27792 12934
rect 27734 12922 27740 12928
rect 27780 12922 27786 12928
rect 24366 12860 24546 12861
rect 28366 12861 28367 13039
rect 28545 12861 28546 13039
rect 32366 13039 32546 13040
rect 31734 12984 31740 12990
rect 31780 12984 31786 12990
rect 31728 12978 31734 12984
rect 31786 12978 31792 12984
rect 31728 12928 31734 12934
rect 31786 12928 31792 12934
rect 31734 12922 31740 12928
rect 31780 12922 31786 12928
rect 28366 12860 28546 12861
rect 32366 12861 32367 13039
rect 32545 12861 32546 13039
rect 36366 13039 36546 13040
rect 35734 12984 35740 12990
rect 35780 12984 35786 12990
rect 35728 12978 35734 12984
rect 35786 12978 35792 12984
rect 35728 12928 35734 12934
rect 35786 12928 35792 12934
rect 35734 12922 35740 12928
rect 35780 12922 35786 12928
rect 32366 12860 32546 12861
rect 36366 12861 36367 13039
rect 36545 12861 36546 13039
rect 39734 12984 39740 12990
rect 39780 12984 39786 12990
rect 39728 12978 39734 12984
rect 39786 12978 39792 12984
rect 39728 12928 39734 12934
rect 39786 12928 39792 12934
rect 39734 12922 39740 12928
rect 39780 12922 39786 12928
rect 36366 12860 36546 12861
rect 3262 12808 3268 12814
rect 3308 12808 3314 12814
rect 7262 12808 7268 12814
rect 7308 12808 7314 12814
rect 11262 12808 11268 12814
rect 11308 12808 11314 12814
rect 15262 12808 15268 12814
rect 15308 12808 15314 12814
rect 19262 12808 19268 12814
rect 19308 12808 19314 12814
rect 23262 12808 23268 12814
rect 23308 12808 23314 12814
rect 27262 12808 27268 12814
rect 27308 12808 27314 12814
rect 31262 12808 31268 12814
rect 31308 12808 31314 12814
rect 35262 12808 35268 12814
rect 35308 12808 35314 12814
rect 39262 12808 39268 12814
rect 39308 12808 39314 12814
rect 3256 12802 3262 12808
rect 3314 12802 3320 12808
rect 7256 12802 7262 12808
rect 7314 12802 7320 12808
rect 11256 12802 11262 12808
rect 11314 12802 11320 12808
rect 15256 12802 15262 12808
rect 15314 12802 15320 12808
rect 19256 12802 19262 12808
rect 19314 12802 19320 12808
rect 23256 12802 23262 12808
rect 23314 12802 23320 12808
rect 27256 12802 27262 12808
rect 27314 12802 27320 12808
rect 31256 12802 31262 12808
rect 31314 12802 31320 12808
rect 35256 12802 35262 12808
rect 35314 12802 35320 12808
rect 39256 12802 39262 12808
rect 39314 12802 39320 12808
rect 3256 12756 3262 12762
rect 3314 12756 3320 12762
rect 7256 12756 7262 12762
rect 7314 12756 7320 12762
rect 11256 12756 11262 12762
rect 11314 12756 11320 12762
rect 15256 12756 15262 12762
rect 15314 12756 15320 12762
rect 19256 12756 19262 12762
rect 19314 12756 19320 12762
rect 23256 12756 23262 12762
rect 23314 12756 23320 12762
rect 27256 12756 27262 12762
rect 27314 12756 27320 12762
rect 31256 12756 31262 12762
rect 31314 12756 31320 12762
rect 35256 12756 35262 12762
rect 35314 12756 35320 12762
rect 39256 12756 39262 12762
rect 39314 12756 39320 12762
rect 3262 12750 3268 12756
rect 3308 12750 3314 12756
rect 7262 12750 7268 12756
rect 7308 12750 7314 12756
rect 11262 12750 11268 12756
rect 11308 12750 11314 12756
rect 15262 12750 15268 12756
rect 15308 12750 15314 12756
rect 19262 12750 19268 12756
rect 19308 12750 19314 12756
rect 23262 12750 23268 12756
rect 23308 12750 23314 12756
rect 27262 12750 27268 12756
rect 27308 12750 27314 12756
rect 31262 12750 31268 12756
rect 31308 12750 31314 12756
rect 35262 12750 35268 12756
rect 35308 12750 35314 12756
rect 39262 12750 39268 12756
rect 39308 12750 39314 12756
rect 2386 12296 2626 12320
rect 2386 12104 2410 12296
rect 2602 12104 2626 12296
rect 2386 12080 2626 12104
rect 6386 12296 6626 12320
rect 6386 12104 6410 12296
rect 6602 12104 6626 12296
rect 6386 12080 6626 12104
rect 10386 12296 10626 12320
rect 10386 12104 10410 12296
rect 10602 12104 10626 12296
rect 10386 12080 10626 12104
rect 14386 12296 14626 12320
rect 14386 12104 14410 12296
rect 14602 12104 14626 12296
rect 14386 12080 14626 12104
rect 18386 12296 18626 12320
rect 18386 12104 18410 12296
rect 18602 12104 18626 12296
rect 18386 12080 18626 12104
rect 22386 12296 22626 12320
rect 22386 12104 22410 12296
rect 22602 12104 22626 12296
rect 22386 12080 22626 12104
rect 26386 12296 26626 12320
rect 26386 12104 26410 12296
rect 26602 12104 26626 12296
rect 26386 12080 26626 12104
rect 30386 12296 30626 12320
rect 30386 12104 30410 12296
rect 30602 12104 30626 12296
rect 30386 12080 30626 12104
rect 34386 12296 34626 12320
rect 34386 12104 34410 12296
rect 34602 12104 34626 12296
rect 34386 12080 34626 12104
rect 38386 12296 38626 12320
rect 38386 12104 38410 12296
rect 38602 12104 38626 12296
rect 38386 12080 38626 12104
rect 1982 11160 2302 11230
rect 366 10916 606 10940
rect 366 10724 390 10916
rect 582 10724 606 10916
rect 1982 10920 2006 11160
rect 2232 10920 2246 11160
rect 2256 10920 2302 11160
rect 5982 11160 6302 11230
rect 1982 10896 2302 10920
rect 4366 10916 4606 10940
rect 366 10700 606 10724
rect 4366 10724 4390 10916
rect 4582 10724 4606 10916
rect 5982 10920 6006 11160
rect 6232 10920 6246 11160
rect 6256 10920 6302 11160
rect 9982 11160 10302 11230
rect 5982 10896 6302 10920
rect 8366 10916 8606 10940
rect 2852 10709 2996 10714
rect 2852 10639 2857 10709
rect 2991 10639 2996 10709
rect 4366 10700 4606 10724
rect 8366 10724 8390 10916
rect 8582 10724 8606 10916
rect 9982 10920 10006 11160
rect 10232 10920 10246 11160
rect 10256 10920 10302 11160
rect 13982 11160 14302 11230
rect 9982 10896 10302 10920
rect 12366 10916 12606 10940
rect 6852 10709 6996 10714
rect 2852 10634 2996 10639
rect 6852 10639 6857 10709
rect 6991 10639 6996 10709
rect 8366 10700 8606 10724
rect 12366 10724 12390 10916
rect 12582 10724 12606 10916
rect 13982 10920 14006 11160
rect 14232 10920 14246 11160
rect 14256 10920 14302 11160
rect 17982 11160 18302 11230
rect 13982 10896 14302 10920
rect 16366 10916 16606 10940
rect 10852 10709 10996 10714
rect 6852 10634 6996 10639
rect 10852 10639 10857 10709
rect 10991 10639 10996 10709
rect 12366 10700 12606 10724
rect 16366 10724 16390 10916
rect 16582 10724 16606 10916
rect 17982 10920 18006 11160
rect 18232 10920 18246 11160
rect 18256 10920 18302 11160
rect 21982 11160 22302 11230
rect 17982 10896 18302 10920
rect 20366 10916 20606 10940
rect 14852 10709 14996 10714
rect 10852 10634 10996 10639
rect 14852 10639 14857 10709
rect 14991 10639 14996 10709
rect 16366 10700 16606 10724
rect 20366 10724 20390 10916
rect 20582 10724 20606 10916
rect 21982 10920 22006 11160
rect 22232 10920 22246 11160
rect 22256 10920 22302 11160
rect 25982 11160 26302 11230
rect 21982 10896 22302 10920
rect 24366 10916 24606 10940
rect 18852 10709 18996 10714
rect 14852 10634 14996 10639
rect 18852 10639 18857 10709
rect 18991 10639 18996 10709
rect 20366 10700 20606 10724
rect 24366 10724 24390 10916
rect 24582 10724 24606 10916
rect 25982 10920 26006 11160
rect 26232 10920 26246 11160
rect 26256 10920 26302 11160
rect 29982 11160 30302 11230
rect 25982 10896 26302 10920
rect 28366 10916 28606 10940
rect 22852 10709 22996 10714
rect 18852 10634 18996 10639
rect 22852 10639 22857 10709
rect 22991 10639 22996 10709
rect 24366 10700 24606 10724
rect 28366 10724 28390 10916
rect 28582 10724 28606 10916
rect 29982 10920 30006 11160
rect 30232 10920 30246 11160
rect 30256 10920 30302 11160
rect 33982 11160 34302 11230
rect 29982 10896 30302 10920
rect 32366 10916 32606 10940
rect 26852 10709 26996 10714
rect 22852 10634 22996 10639
rect 26852 10639 26857 10709
rect 26991 10639 26996 10709
rect 28366 10700 28606 10724
rect 32366 10724 32390 10916
rect 32582 10724 32606 10916
rect 33982 10920 34006 11160
rect 34232 10920 34246 11160
rect 34256 10920 34302 11160
rect 37982 11160 38302 11230
rect 33982 10896 34302 10920
rect 36366 10916 36606 10940
rect 30852 10709 30996 10714
rect 26852 10634 26996 10639
rect 30852 10639 30857 10709
rect 30991 10639 30996 10709
rect 32366 10700 32606 10724
rect 36366 10724 36390 10916
rect 36582 10724 36606 10916
rect 37982 10920 38006 11160
rect 38232 10920 38246 11160
rect 38256 10920 38302 11160
rect 37982 10896 38302 10920
rect 34852 10709 34996 10714
rect 30852 10634 30996 10639
rect 34852 10639 34857 10709
rect 34991 10639 34996 10709
rect 36366 10700 36606 10724
rect 38852 10709 38996 10714
rect 34852 10634 34996 10639
rect 38852 10639 38857 10709
rect 38991 10639 38996 10709
rect 38852 10634 38996 10639
rect 2366 10559 2546 10560
rect 2366 10381 2367 10559
rect 2545 10381 2546 10559
rect 2366 10380 2546 10381
rect 6366 10559 6546 10560
rect 6366 10381 6367 10559
rect 6545 10381 6546 10559
rect 6366 10380 6546 10381
rect 10366 10559 10546 10560
rect 10366 10381 10367 10559
rect 10545 10381 10546 10559
rect 10366 10380 10546 10381
rect 14366 10559 14546 10560
rect 14366 10381 14367 10559
rect 14545 10381 14546 10559
rect 14366 10380 14546 10381
rect 18366 10559 18546 10560
rect 18366 10381 18367 10559
rect 18545 10381 18546 10559
rect 18366 10380 18546 10381
rect 22366 10559 22546 10560
rect 22366 10381 22367 10559
rect 22545 10381 22546 10559
rect 22366 10380 22546 10381
rect 26366 10559 26546 10560
rect 26366 10381 26367 10559
rect 26545 10381 26546 10559
rect 26366 10380 26546 10381
rect 30366 10559 30546 10560
rect 30366 10381 30367 10559
rect 30545 10381 30546 10559
rect 30366 10380 30546 10381
rect 34366 10559 34546 10560
rect 34366 10381 34367 10559
rect 34545 10381 34546 10559
rect 34366 10380 34546 10381
rect 38366 10559 38546 10560
rect 38366 10381 38367 10559
rect 38545 10381 38546 10559
rect 38366 10380 38546 10381
rect 366 10039 546 10040
rect 366 9861 367 10039
rect 545 9861 546 10039
rect 4366 10039 4546 10040
rect 3734 9984 3740 9990
rect 3780 9984 3786 9990
rect 3728 9978 3734 9984
rect 3786 9978 3792 9984
rect 3728 9928 3734 9934
rect 3786 9928 3792 9934
rect 3734 9922 3740 9928
rect 3780 9922 3786 9928
rect 366 9860 546 9861
rect 4366 9861 4367 10039
rect 4545 9861 4546 10039
rect 8366 10039 8546 10040
rect 7734 9984 7740 9990
rect 7780 9984 7786 9990
rect 7728 9978 7734 9984
rect 7786 9978 7792 9984
rect 7728 9928 7734 9934
rect 7786 9928 7792 9934
rect 7734 9922 7740 9928
rect 7780 9922 7786 9928
rect 4366 9860 4546 9861
rect 8366 9861 8367 10039
rect 8545 9861 8546 10039
rect 12366 10039 12546 10040
rect 11734 9984 11740 9990
rect 11780 9984 11786 9990
rect 11728 9978 11734 9984
rect 11786 9978 11792 9984
rect 11728 9928 11734 9934
rect 11786 9928 11792 9934
rect 11734 9922 11740 9928
rect 11780 9922 11786 9928
rect 8366 9860 8546 9861
rect 12366 9861 12367 10039
rect 12545 9861 12546 10039
rect 16366 10039 16546 10040
rect 15734 9984 15740 9990
rect 15780 9984 15786 9990
rect 15728 9978 15734 9984
rect 15786 9978 15792 9984
rect 15728 9928 15734 9934
rect 15786 9928 15792 9934
rect 15734 9922 15740 9928
rect 15780 9922 15786 9928
rect 12366 9860 12546 9861
rect 16366 9861 16367 10039
rect 16545 9861 16546 10039
rect 20366 10039 20546 10040
rect 19734 9984 19740 9990
rect 19780 9984 19786 9990
rect 19728 9978 19734 9984
rect 19786 9978 19792 9984
rect 19728 9928 19734 9934
rect 19786 9928 19792 9934
rect 19734 9922 19740 9928
rect 19780 9922 19786 9928
rect 16366 9860 16546 9861
rect 20366 9861 20367 10039
rect 20545 9861 20546 10039
rect 24366 10039 24546 10040
rect 23734 9984 23740 9990
rect 23780 9984 23786 9990
rect 23728 9978 23734 9984
rect 23786 9978 23792 9984
rect 23728 9928 23734 9934
rect 23786 9928 23792 9934
rect 23734 9922 23740 9928
rect 23780 9922 23786 9928
rect 20366 9860 20546 9861
rect 24366 9861 24367 10039
rect 24545 9861 24546 10039
rect 28366 10039 28546 10040
rect 27734 9984 27740 9990
rect 27780 9984 27786 9990
rect 27728 9978 27734 9984
rect 27786 9978 27792 9984
rect 27728 9928 27734 9934
rect 27786 9928 27792 9934
rect 27734 9922 27740 9928
rect 27780 9922 27786 9928
rect 24366 9860 24546 9861
rect 28366 9861 28367 10039
rect 28545 9861 28546 10039
rect 32366 10039 32546 10040
rect 31734 9984 31740 9990
rect 31780 9984 31786 9990
rect 31728 9978 31734 9984
rect 31786 9978 31792 9984
rect 31728 9928 31734 9934
rect 31786 9928 31792 9934
rect 31734 9922 31740 9928
rect 31780 9922 31786 9928
rect 28366 9860 28546 9861
rect 32366 9861 32367 10039
rect 32545 9861 32546 10039
rect 36366 10039 36546 10040
rect 35734 9984 35740 9990
rect 35780 9984 35786 9990
rect 35728 9978 35734 9984
rect 35786 9978 35792 9984
rect 35728 9928 35734 9934
rect 35786 9928 35792 9934
rect 35734 9922 35740 9928
rect 35780 9922 35786 9928
rect 32366 9860 32546 9861
rect 36366 9861 36367 10039
rect 36545 9861 36546 10039
rect 39734 9984 39740 9990
rect 39780 9984 39786 9990
rect 39728 9978 39734 9984
rect 39786 9978 39792 9984
rect 39728 9928 39734 9934
rect 39786 9928 39792 9934
rect 39734 9922 39740 9928
rect 39780 9922 39786 9928
rect 36366 9860 36546 9861
rect 3262 9808 3268 9814
rect 3308 9808 3314 9814
rect 7262 9808 7268 9814
rect 7308 9808 7314 9814
rect 11262 9808 11268 9814
rect 11308 9808 11314 9814
rect 15262 9808 15268 9814
rect 15308 9808 15314 9814
rect 19262 9808 19268 9814
rect 19308 9808 19314 9814
rect 23262 9808 23268 9814
rect 23308 9808 23314 9814
rect 27262 9808 27268 9814
rect 27308 9808 27314 9814
rect 31262 9808 31268 9814
rect 31308 9808 31314 9814
rect 35262 9808 35268 9814
rect 35308 9808 35314 9814
rect 39262 9808 39268 9814
rect 39308 9808 39314 9814
rect 3256 9802 3262 9808
rect 3314 9802 3320 9808
rect 7256 9802 7262 9808
rect 7314 9802 7320 9808
rect 11256 9802 11262 9808
rect 11314 9802 11320 9808
rect 15256 9802 15262 9808
rect 15314 9802 15320 9808
rect 19256 9802 19262 9808
rect 19314 9802 19320 9808
rect 23256 9802 23262 9808
rect 23314 9802 23320 9808
rect 27256 9802 27262 9808
rect 27314 9802 27320 9808
rect 31256 9802 31262 9808
rect 31314 9802 31320 9808
rect 35256 9802 35262 9808
rect 35314 9802 35320 9808
rect 39256 9802 39262 9808
rect 39314 9802 39320 9808
rect 3256 9756 3262 9762
rect 3314 9756 3320 9762
rect 7256 9756 7262 9762
rect 7314 9756 7320 9762
rect 11256 9756 11262 9762
rect 11314 9756 11320 9762
rect 15256 9756 15262 9762
rect 15314 9756 15320 9762
rect 19256 9756 19262 9762
rect 19314 9756 19320 9762
rect 23256 9756 23262 9762
rect 23314 9756 23320 9762
rect 27256 9756 27262 9762
rect 27314 9756 27320 9762
rect 31256 9756 31262 9762
rect 31314 9756 31320 9762
rect 35256 9756 35262 9762
rect 35314 9756 35320 9762
rect 39256 9756 39262 9762
rect 39314 9756 39320 9762
rect 3262 9750 3268 9756
rect 3308 9750 3314 9756
rect 7262 9750 7268 9756
rect 7308 9750 7314 9756
rect 11262 9750 11268 9756
rect 11308 9750 11314 9756
rect 15262 9750 15268 9756
rect 15308 9750 15314 9756
rect 19262 9750 19268 9756
rect 19308 9750 19314 9756
rect 23262 9750 23268 9756
rect 23308 9750 23314 9756
rect 27262 9750 27268 9756
rect 27308 9750 27314 9756
rect 31262 9750 31268 9756
rect 31308 9750 31314 9756
rect 35262 9750 35268 9756
rect 35308 9750 35314 9756
rect 39262 9750 39268 9756
rect 39308 9750 39314 9756
rect 2386 9296 2626 9320
rect 2386 9104 2410 9296
rect 2602 9104 2626 9296
rect 2386 9080 2626 9104
rect 6386 9296 6626 9320
rect 6386 9104 6410 9296
rect 6602 9104 6626 9296
rect 6386 9080 6626 9104
rect 10386 9296 10626 9320
rect 10386 9104 10410 9296
rect 10602 9104 10626 9296
rect 10386 9080 10626 9104
rect 14386 9296 14626 9320
rect 14386 9104 14410 9296
rect 14602 9104 14626 9296
rect 14386 9080 14626 9104
rect 18386 9296 18626 9320
rect 18386 9104 18410 9296
rect 18602 9104 18626 9296
rect 18386 9080 18626 9104
rect 22386 9296 22626 9320
rect 22386 9104 22410 9296
rect 22602 9104 22626 9296
rect 22386 9080 22626 9104
rect 26386 9296 26626 9320
rect 26386 9104 26410 9296
rect 26602 9104 26626 9296
rect 26386 9080 26626 9104
rect 30386 9296 30626 9320
rect 30386 9104 30410 9296
rect 30602 9104 30626 9296
rect 30386 9080 30626 9104
rect 34386 9296 34626 9320
rect 34386 9104 34410 9296
rect 34602 9104 34626 9296
rect 34386 9080 34626 9104
rect 38386 9296 38626 9320
rect 38386 9104 38410 9296
rect 38602 9104 38626 9296
rect 38386 9080 38626 9104
rect 1982 8160 2302 8230
rect 366 7916 606 7940
rect 366 7724 390 7916
rect 582 7724 606 7916
rect 1982 7920 2006 8160
rect 2232 7920 2246 8160
rect 2256 7920 2302 8160
rect 5982 8160 6302 8230
rect 1982 7896 2302 7920
rect 4366 7916 4606 7940
rect 366 7700 606 7724
rect 4366 7724 4390 7916
rect 4582 7724 4606 7916
rect 5982 7920 6006 8160
rect 6232 7920 6246 8160
rect 6256 7920 6302 8160
rect 9982 8160 10302 8230
rect 5982 7896 6302 7920
rect 8366 7916 8606 7940
rect 2852 7709 2996 7714
rect 2852 7639 2857 7709
rect 2991 7639 2996 7709
rect 4366 7700 4606 7724
rect 8366 7724 8390 7916
rect 8582 7724 8606 7916
rect 9982 7920 10006 8160
rect 10232 7920 10246 8160
rect 10256 7920 10302 8160
rect 13982 8160 14302 8230
rect 9982 7896 10302 7920
rect 12366 7916 12606 7940
rect 6852 7709 6996 7714
rect 2852 7634 2996 7639
rect 6852 7639 6857 7709
rect 6991 7639 6996 7709
rect 8366 7700 8606 7724
rect 12366 7724 12390 7916
rect 12582 7724 12606 7916
rect 13982 7920 14006 8160
rect 14232 7920 14246 8160
rect 14256 7920 14302 8160
rect 17982 8160 18302 8230
rect 13982 7896 14302 7920
rect 16366 7916 16606 7940
rect 10852 7709 10996 7714
rect 6852 7634 6996 7639
rect 10852 7639 10857 7709
rect 10991 7639 10996 7709
rect 12366 7700 12606 7724
rect 16366 7724 16390 7916
rect 16582 7724 16606 7916
rect 17982 7920 18006 8160
rect 18232 7920 18246 8160
rect 18256 7920 18302 8160
rect 21982 8160 22302 8230
rect 17982 7896 18302 7920
rect 20366 7916 20606 7940
rect 14852 7709 14996 7714
rect 10852 7634 10996 7639
rect 14852 7639 14857 7709
rect 14991 7639 14996 7709
rect 16366 7700 16606 7724
rect 20366 7724 20390 7916
rect 20582 7724 20606 7916
rect 21982 7920 22006 8160
rect 22232 7920 22246 8160
rect 22256 7920 22302 8160
rect 25982 8160 26302 8230
rect 21982 7896 22302 7920
rect 24366 7916 24606 7940
rect 18852 7709 18996 7714
rect 14852 7634 14996 7639
rect 18852 7639 18857 7709
rect 18991 7639 18996 7709
rect 20366 7700 20606 7724
rect 24366 7724 24390 7916
rect 24582 7724 24606 7916
rect 25982 7920 26006 8160
rect 26232 7920 26246 8160
rect 26256 7920 26302 8160
rect 29982 8160 30302 8230
rect 25982 7896 26302 7920
rect 28366 7916 28606 7940
rect 22852 7709 22996 7714
rect 18852 7634 18996 7639
rect 22852 7639 22857 7709
rect 22991 7639 22996 7709
rect 24366 7700 24606 7724
rect 28366 7724 28390 7916
rect 28582 7724 28606 7916
rect 29982 7920 30006 8160
rect 30232 7920 30246 8160
rect 30256 7920 30302 8160
rect 33982 8160 34302 8230
rect 29982 7896 30302 7920
rect 32366 7916 32606 7940
rect 26852 7709 26996 7714
rect 22852 7634 22996 7639
rect 26852 7639 26857 7709
rect 26991 7639 26996 7709
rect 28366 7700 28606 7724
rect 32366 7724 32390 7916
rect 32582 7724 32606 7916
rect 33982 7920 34006 8160
rect 34232 7920 34246 8160
rect 34256 7920 34302 8160
rect 37982 8160 38302 8230
rect 33982 7896 34302 7920
rect 36366 7916 36606 7940
rect 30852 7709 30996 7714
rect 26852 7634 26996 7639
rect 30852 7639 30857 7709
rect 30991 7639 30996 7709
rect 32366 7700 32606 7724
rect 36366 7724 36390 7916
rect 36582 7724 36606 7916
rect 37982 7920 38006 8160
rect 38232 7920 38246 8160
rect 38256 7920 38302 8160
rect 37982 7896 38302 7920
rect 34852 7709 34996 7714
rect 30852 7634 30996 7639
rect 34852 7639 34857 7709
rect 34991 7639 34996 7709
rect 36366 7700 36606 7724
rect 38852 7709 38996 7714
rect 34852 7634 34996 7639
rect 38852 7639 38857 7709
rect 38991 7639 38996 7709
rect 38852 7634 38996 7639
rect 2366 7559 2546 7560
rect 2366 7381 2367 7559
rect 2545 7381 2546 7559
rect 2366 7380 2546 7381
rect 6366 7559 6546 7560
rect 6366 7381 6367 7559
rect 6545 7381 6546 7559
rect 6366 7380 6546 7381
rect 10366 7559 10546 7560
rect 10366 7381 10367 7559
rect 10545 7381 10546 7559
rect 10366 7380 10546 7381
rect 14366 7559 14546 7560
rect 14366 7381 14367 7559
rect 14545 7381 14546 7559
rect 14366 7380 14546 7381
rect 18366 7559 18546 7560
rect 18366 7381 18367 7559
rect 18545 7381 18546 7559
rect 18366 7380 18546 7381
rect 22366 7559 22546 7560
rect 22366 7381 22367 7559
rect 22545 7381 22546 7559
rect 22366 7380 22546 7381
rect 26366 7559 26546 7560
rect 26366 7381 26367 7559
rect 26545 7381 26546 7559
rect 26366 7380 26546 7381
rect 30366 7559 30546 7560
rect 30366 7381 30367 7559
rect 30545 7381 30546 7559
rect 30366 7380 30546 7381
rect 34366 7559 34546 7560
rect 34366 7381 34367 7559
rect 34545 7381 34546 7559
rect 34366 7380 34546 7381
rect 38366 7559 38546 7560
rect 38366 7381 38367 7559
rect 38545 7381 38546 7559
rect 38366 7380 38546 7381
rect 366 7039 546 7040
rect 366 6861 367 7039
rect 545 6861 546 7039
rect 4366 7039 4546 7040
rect 3734 6984 3740 6990
rect 3780 6984 3786 6990
rect 3728 6978 3734 6984
rect 3786 6978 3792 6984
rect 3728 6928 3734 6934
rect 3786 6928 3792 6934
rect 3734 6922 3740 6928
rect 3780 6922 3786 6928
rect 366 6860 546 6861
rect 4366 6861 4367 7039
rect 4545 6861 4546 7039
rect 8366 7039 8546 7040
rect 7734 6984 7740 6990
rect 7780 6984 7786 6990
rect 7728 6978 7734 6984
rect 7786 6978 7792 6984
rect 7728 6928 7734 6934
rect 7786 6928 7792 6934
rect 7734 6922 7740 6928
rect 7780 6922 7786 6928
rect 4366 6860 4546 6861
rect 8366 6861 8367 7039
rect 8545 6861 8546 7039
rect 12366 7039 12546 7040
rect 11734 6984 11740 6990
rect 11780 6984 11786 6990
rect 11728 6978 11734 6984
rect 11786 6978 11792 6984
rect 11728 6928 11734 6934
rect 11786 6928 11792 6934
rect 11734 6922 11740 6928
rect 11780 6922 11786 6928
rect 8366 6860 8546 6861
rect 12366 6861 12367 7039
rect 12545 6861 12546 7039
rect 16366 7039 16546 7040
rect 15734 6984 15740 6990
rect 15780 6984 15786 6990
rect 15728 6978 15734 6984
rect 15786 6978 15792 6984
rect 15728 6928 15734 6934
rect 15786 6928 15792 6934
rect 15734 6922 15740 6928
rect 15780 6922 15786 6928
rect 12366 6860 12546 6861
rect 16366 6861 16367 7039
rect 16545 6861 16546 7039
rect 20366 7039 20546 7040
rect 19734 6984 19740 6990
rect 19780 6984 19786 6990
rect 19728 6978 19734 6984
rect 19786 6978 19792 6984
rect 19728 6928 19734 6934
rect 19786 6928 19792 6934
rect 19734 6922 19740 6928
rect 19780 6922 19786 6928
rect 16366 6860 16546 6861
rect 20366 6861 20367 7039
rect 20545 6861 20546 7039
rect 24366 7039 24546 7040
rect 23734 6984 23740 6990
rect 23780 6984 23786 6990
rect 23728 6978 23734 6984
rect 23786 6978 23792 6984
rect 23728 6928 23734 6934
rect 23786 6928 23792 6934
rect 23734 6922 23740 6928
rect 23780 6922 23786 6928
rect 20366 6860 20546 6861
rect 24366 6861 24367 7039
rect 24545 6861 24546 7039
rect 28366 7039 28546 7040
rect 27734 6984 27740 6990
rect 27780 6984 27786 6990
rect 27728 6978 27734 6984
rect 27786 6978 27792 6984
rect 27728 6928 27734 6934
rect 27786 6928 27792 6934
rect 27734 6922 27740 6928
rect 27780 6922 27786 6928
rect 24366 6860 24546 6861
rect 28366 6861 28367 7039
rect 28545 6861 28546 7039
rect 32366 7039 32546 7040
rect 31734 6984 31740 6990
rect 31780 6984 31786 6990
rect 31728 6978 31734 6984
rect 31786 6978 31792 6984
rect 31728 6928 31734 6934
rect 31786 6928 31792 6934
rect 31734 6922 31740 6928
rect 31780 6922 31786 6928
rect 28366 6860 28546 6861
rect 32366 6861 32367 7039
rect 32545 6861 32546 7039
rect 36366 7039 36546 7040
rect 35734 6984 35740 6990
rect 35780 6984 35786 6990
rect 35728 6978 35734 6984
rect 35786 6978 35792 6984
rect 35728 6928 35734 6934
rect 35786 6928 35792 6934
rect 35734 6922 35740 6928
rect 35780 6922 35786 6928
rect 32366 6860 32546 6861
rect 36366 6861 36367 7039
rect 36545 6861 36546 7039
rect 39734 6984 39740 6990
rect 39780 6984 39786 6990
rect 39728 6978 39734 6984
rect 39786 6978 39792 6984
rect 39728 6928 39734 6934
rect 39786 6928 39792 6934
rect 39734 6922 39740 6928
rect 39780 6922 39786 6928
rect 36366 6860 36546 6861
rect 3262 6808 3268 6814
rect 3308 6808 3314 6814
rect 7262 6808 7268 6814
rect 7308 6808 7314 6814
rect 11262 6808 11268 6814
rect 11308 6808 11314 6814
rect 15262 6808 15268 6814
rect 15308 6808 15314 6814
rect 19262 6808 19268 6814
rect 19308 6808 19314 6814
rect 23262 6808 23268 6814
rect 23308 6808 23314 6814
rect 27262 6808 27268 6814
rect 27308 6808 27314 6814
rect 31262 6808 31268 6814
rect 31308 6808 31314 6814
rect 35262 6808 35268 6814
rect 35308 6808 35314 6814
rect 39262 6808 39268 6814
rect 39308 6808 39314 6814
rect 3256 6802 3262 6808
rect 3314 6802 3320 6808
rect 7256 6802 7262 6808
rect 7314 6802 7320 6808
rect 11256 6802 11262 6808
rect 11314 6802 11320 6808
rect 15256 6802 15262 6808
rect 15314 6802 15320 6808
rect 19256 6802 19262 6808
rect 19314 6802 19320 6808
rect 23256 6802 23262 6808
rect 23314 6802 23320 6808
rect 27256 6802 27262 6808
rect 27314 6802 27320 6808
rect 31256 6802 31262 6808
rect 31314 6802 31320 6808
rect 35256 6802 35262 6808
rect 35314 6802 35320 6808
rect 39256 6802 39262 6808
rect 39314 6802 39320 6808
rect 3256 6756 3262 6762
rect 3314 6756 3320 6762
rect 7256 6756 7262 6762
rect 7314 6756 7320 6762
rect 11256 6756 11262 6762
rect 11314 6756 11320 6762
rect 15256 6756 15262 6762
rect 15314 6756 15320 6762
rect 19256 6756 19262 6762
rect 19314 6756 19320 6762
rect 23256 6756 23262 6762
rect 23314 6756 23320 6762
rect 27256 6756 27262 6762
rect 27314 6756 27320 6762
rect 31256 6756 31262 6762
rect 31314 6756 31320 6762
rect 35256 6756 35262 6762
rect 35314 6756 35320 6762
rect 39256 6756 39262 6762
rect 39314 6756 39320 6762
rect 3262 6750 3268 6756
rect 3308 6750 3314 6756
rect 7262 6750 7268 6756
rect 7308 6750 7314 6756
rect 11262 6750 11268 6756
rect 11308 6750 11314 6756
rect 15262 6750 15268 6756
rect 15308 6750 15314 6756
rect 19262 6750 19268 6756
rect 19308 6750 19314 6756
rect 23262 6750 23268 6756
rect 23308 6750 23314 6756
rect 27262 6750 27268 6756
rect 27308 6750 27314 6756
rect 31262 6750 31268 6756
rect 31308 6750 31314 6756
rect 35262 6750 35268 6756
rect 35308 6750 35314 6756
rect 39262 6750 39268 6756
rect 39308 6750 39314 6756
rect 2386 6296 2626 6320
rect 2386 6104 2410 6296
rect 2602 6104 2626 6296
rect 2386 6080 2626 6104
rect 6386 6296 6626 6320
rect 6386 6104 6410 6296
rect 6602 6104 6626 6296
rect 6386 6080 6626 6104
rect 10386 6296 10626 6320
rect 10386 6104 10410 6296
rect 10602 6104 10626 6296
rect 10386 6080 10626 6104
rect 14386 6296 14626 6320
rect 14386 6104 14410 6296
rect 14602 6104 14626 6296
rect 14386 6080 14626 6104
rect 18386 6296 18626 6320
rect 18386 6104 18410 6296
rect 18602 6104 18626 6296
rect 18386 6080 18626 6104
rect 22386 6296 22626 6320
rect 22386 6104 22410 6296
rect 22602 6104 22626 6296
rect 22386 6080 22626 6104
rect 26386 6296 26626 6320
rect 26386 6104 26410 6296
rect 26602 6104 26626 6296
rect 26386 6080 26626 6104
rect 30386 6296 30626 6320
rect 30386 6104 30410 6296
rect 30602 6104 30626 6296
rect 30386 6080 30626 6104
rect 34386 6296 34626 6320
rect 34386 6104 34410 6296
rect 34602 6104 34626 6296
rect 34386 6080 34626 6104
rect 38386 6296 38626 6320
rect 38386 6104 38410 6296
rect 38602 6104 38626 6296
rect 38386 6080 38626 6104
rect 1982 5160 2302 5230
rect 366 4916 606 4940
rect 366 4724 390 4916
rect 582 4724 606 4916
rect 1982 4920 2006 5160
rect 2232 4920 2246 5160
rect 2256 4920 2302 5160
rect 5982 5160 6302 5230
rect 1982 4896 2302 4920
rect 4366 4916 4606 4940
rect 366 4700 606 4724
rect 4366 4724 4390 4916
rect 4582 4724 4606 4916
rect 5982 4920 6006 5160
rect 6232 4920 6246 5160
rect 6256 4920 6302 5160
rect 9982 5160 10302 5230
rect 5982 4896 6302 4920
rect 8366 4916 8606 4940
rect 2852 4709 2996 4714
rect 2852 4639 2857 4709
rect 2991 4639 2996 4709
rect 4366 4700 4606 4724
rect 8366 4724 8390 4916
rect 8582 4724 8606 4916
rect 9982 4920 10006 5160
rect 10232 4920 10246 5160
rect 10256 4920 10302 5160
rect 13982 5160 14302 5230
rect 9982 4896 10302 4920
rect 12366 4916 12606 4940
rect 6852 4709 6996 4714
rect 2852 4634 2996 4639
rect 6852 4639 6857 4709
rect 6991 4639 6996 4709
rect 8366 4700 8606 4724
rect 12366 4724 12390 4916
rect 12582 4724 12606 4916
rect 13982 4920 14006 5160
rect 14232 4920 14246 5160
rect 14256 4920 14302 5160
rect 17982 5160 18302 5230
rect 13982 4896 14302 4920
rect 16366 4916 16606 4940
rect 10852 4709 10996 4714
rect 6852 4634 6996 4639
rect 10852 4639 10857 4709
rect 10991 4639 10996 4709
rect 12366 4700 12606 4724
rect 16366 4724 16390 4916
rect 16582 4724 16606 4916
rect 17982 4920 18006 5160
rect 18232 4920 18246 5160
rect 18256 4920 18302 5160
rect 21982 5160 22302 5230
rect 17982 4896 18302 4920
rect 20366 4916 20606 4940
rect 14852 4709 14996 4714
rect 10852 4634 10996 4639
rect 14852 4639 14857 4709
rect 14991 4639 14996 4709
rect 16366 4700 16606 4724
rect 20366 4724 20390 4916
rect 20582 4724 20606 4916
rect 21982 4920 22006 5160
rect 22232 4920 22246 5160
rect 22256 4920 22302 5160
rect 25982 5160 26302 5230
rect 21982 4896 22302 4920
rect 24366 4916 24606 4940
rect 18852 4709 18996 4714
rect 14852 4634 14996 4639
rect 18852 4639 18857 4709
rect 18991 4639 18996 4709
rect 20366 4700 20606 4724
rect 24366 4724 24390 4916
rect 24582 4724 24606 4916
rect 25982 4920 26006 5160
rect 26232 4920 26246 5160
rect 26256 4920 26302 5160
rect 29982 5160 30302 5230
rect 25982 4896 26302 4920
rect 28366 4916 28606 4940
rect 22852 4709 22996 4714
rect 18852 4634 18996 4639
rect 22852 4639 22857 4709
rect 22991 4639 22996 4709
rect 24366 4700 24606 4724
rect 28366 4724 28390 4916
rect 28582 4724 28606 4916
rect 29982 4920 30006 5160
rect 30232 4920 30246 5160
rect 30256 4920 30302 5160
rect 33982 5160 34302 5230
rect 29982 4896 30302 4920
rect 32366 4916 32606 4940
rect 26852 4709 26996 4714
rect 22852 4634 22996 4639
rect 26852 4639 26857 4709
rect 26991 4639 26996 4709
rect 28366 4700 28606 4724
rect 32366 4724 32390 4916
rect 32582 4724 32606 4916
rect 33982 4920 34006 5160
rect 34232 4920 34246 5160
rect 34256 4920 34302 5160
rect 37982 5160 38302 5230
rect 33982 4896 34302 4920
rect 36366 4916 36606 4940
rect 30852 4709 30996 4714
rect 26852 4634 26996 4639
rect 30852 4639 30857 4709
rect 30991 4639 30996 4709
rect 32366 4700 32606 4724
rect 36366 4724 36390 4916
rect 36582 4724 36606 4916
rect 37982 4920 38006 5160
rect 38232 4920 38246 5160
rect 38256 4920 38302 5160
rect 37982 4896 38302 4920
rect 34852 4709 34996 4714
rect 30852 4634 30996 4639
rect 34852 4639 34857 4709
rect 34991 4639 34996 4709
rect 36366 4700 36606 4724
rect 38852 4709 38996 4714
rect 34852 4634 34996 4639
rect 38852 4639 38857 4709
rect 38991 4639 38996 4709
rect 38852 4634 38996 4639
rect 2366 4559 2546 4560
rect 2366 4381 2367 4559
rect 2545 4381 2546 4559
rect 2366 4380 2546 4381
rect 6366 4559 6546 4560
rect 6366 4381 6367 4559
rect 6545 4381 6546 4559
rect 6366 4380 6546 4381
rect 10366 4559 10546 4560
rect 10366 4381 10367 4559
rect 10545 4381 10546 4559
rect 10366 4380 10546 4381
rect 14366 4559 14546 4560
rect 14366 4381 14367 4559
rect 14545 4381 14546 4559
rect 14366 4380 14546 4381
rect 18366 4559 18546 4560
rect 18366 4381 18367 4559
rect 18545 4381 18546 4559
rect 18366 4380 18546 4381
rect 22366 4559 22546 4560
rect 22366 4381 22367 4559
rect 22545 4381 22546 4559
rect 22366 4380 22546 4381
rect 26366 4559 26546 4560
rect 26366 4381 26367 4559
rect 26545 4381 26546 4559
rect 26366 4380 26546 4381
rect 30366 4559 30546 4560
rect 30366 4381 30367 4559
rect 30545 4381 30546 4559
rect 30366 4380 30546 4381
rect 34366 4559 34546 4560
rect 34366 4381 34367 4559
rect 34545 4381 34546 4559
rect 34366 4380 34546 4381
rect 38366 4559 38546 4560
rect 38366 4381 38367 4559
rect 38545 4381 38546 4559
rect 38366 4380 38546 4381
rect 366 4039 546 4040
rect 366 3861 367 4039
rect 545 3861 546 4039
rect 4366 4039 4546 4040
rect 3734 3984 3740 3990
rect 3780 3984 3786 3990
rect 3728 3978 3734 3984
rect 3786 3978 3792 3984
rect 3728 3928 3734 3934
rect 3786 3928 3792 3934
rect 3734 3922 3740 3928
rect 3780 3922 3786 3928
rect 366 3860 546 3861
rect 4366 3861 4367 4039
rect 4545 3861 4546 4039
rect 8366 4039 8546 4040
rect 7734 3984 7740 3990
rect 7780 3984 7786 3990
rect 7728 3978 7734 3984
rect 7786 3978 7792 3984
rect 7728 3928 7734 3934
rect 7786 3928 7792 3934
rect 7734 3922 7740 3928
rect 7780 3922 7786 3928
rect 4366 3860 4546 3861
rect 8366 3861 8367 4039
rect 8545 3861 8546 4039
rect 12366 4039 12546 4040
rect 11734 3984 11740 3990
rect 11780 3984 11786 3990
rect 11728 3978 11734 3984
rect 11786 3978 11792 3984
rect 11728 3928 11734 3934
rect 11786 3928 11792 3934
rect 11734 3922 11740 3928
rect 11780 3922 11786 3928
rect 8366 3860 8546 3861
rect 12366 3861 12367 4039
rect 12545 3861 12546 4039
rect 16366 4039 16546 4040
rect 15734 3984 15740 3990
rect 15780 3984 15786 3990
rect 15728 3978 15734 3984
rect 15786 3978 15792 3984
rect 15728 3928 15734 3934
rect 15786 3928 15792 3934
rect 15734 3922 15740 3928
rect 15780 3922 15786 3928
rect 12366 3860 12546 3861
rect 16366 3861 16367 4039
rect 16545 3861 16546 4039
rect 20366 4039 20546 4040
rect 19734 3984 19740 3990
rect 19780 3984 19786 3990
rect 19728 3978 19734 3984
rect 19786 3978 19792 3984
rect 19728 3928 19734 3934
rect 19786 3928 19792 3934
rect 19734 3922 19740 3928
rect 19780 3922 19786 3928
rect 16366 3860 16546 3861
rect 20366 3861 20367 4039
rect 20545 3861 20546 4039
rect 24366 4039 24546 4040
rect 23734 3984 23740 3990
rect 23780 3984 23786 3990
rect 23728 3978 23734 3984
rect 23786 3978 23792 3984
rect 23728 3928 23734 3934
rect 23786 3928 23792 3934
rect 23734 3922 23740 3928
rect 23780 3922 23786 3928
rect 20366 3860 20546 3861
rect 24366 3861 24367 4039
rect 24545 3861 24546 4039
rect 28366 4039 28546 4040
rect 27734 3984 27740 3990
rect 27780 3984 27786 3990
rect 27728 3978 27734 3984
rect 27786 3978 27792 3984
rect 27728 3928 27734 3934
rect 27786 3928 27792 3934
rect 27734 3922 27740 3928
rect 27780 3922 27786 3928
rect 24366 3860 24546 3861
rect 28366 3861 28367 4039
rect 28545 3861 28546 4039
rect 32366 4039 32546 4040
rect 31734 3984 31740 3990
rect 31780 3984 31786 3990
rect 31728 3978 31734 3984
rect 31786 3978 31792 3984
rect 31728 3928 31734 3934
rect 31786 3928 31792 3934
rect 31734 3922 31740 3928
rect 31780 3922 31786 3928
rect 28366 3860 28546 3861
rect 32366 3861 32367 4039
rect 32545 3861 32546 4039
rect 36366 4039 36546 4040
rect 35734 3984 35740 3990
rect 35780 3984 35786 3990
rect 35728 3978 35734 3984
rect 35786 3978 35792 3984
rect 35728 3928 35734 3934
rect 35786 3928 35792 3934
rect 35734 3922 35740 3928
rect 35780 3922 35786 3928
rect 32366 3860 32546 3861
rect 36366 3861 36367 4039
rect 36545 3861 36546 4039
rect 39734 3984 39740 3990
rect 39780 3984 39786 3990
rect 39728 3978 39734 3984
rect 39786 3978 39792 3984
rect 39728 3928 39734 3934
rect 39786 3928 39792 3934
rect 39734 3922 39740 3928
rect 39780 3922 39786 3928
rect 36366 3860 36546 3861
rect 3262 3808 3268 3814
rect 3308 3808 3314 3814
rect 7262 3808 7268 3814
rect 7308 3808 7314 3814
rect 11262 3808 11268 3814
rect 11308 3808 11314 3814
rect 15262 3808 15268 3814
rect 15308 3808 15314 3814
rect 19262 3808 19268 3814
rect 19308 3808 19314 3814
rect 23262 3808 23268 3814
rect 23308 3808 23314 3814
rect 27262 3808 27268 3814
rect 27308 3808 27314 3814
rect 31262 3808 31268 3814
rect 31308 3808 31314 3814
rect 35262 3808 35268 3814
rect 35308 3808 35314 3814
rect 39262 3808 39268 3814
rect 39308 3808 39314 3814
rect 3256 3802 3262 3808
rect 3314 3802 3320 3808
rect 7256 3802 7262 3808
rect 7314 3802 7320 3808
rect 11256 3802 11262 3808
rect 11314 3802 11320 3808
rect 15256 3802 15262 3808
rect 15314 3802 15320 3808
rect 19256 3802 19262 3808
rect 19314 3802 19320 3808
rect 23256 3802 23262 3808
rect 23314 3802 23320 3808
rect 27256 3802 27262 3808
rect 27314 3802 27320 3808
rect 31256 3802 31262 3808
rect 31314 3802 31320 3808
rect 35256 3802 35262 3808
rect 35314 3802 35320 3808
rect 39256 3802 39262 3808
rect 39314 3802 39320 3808
rect 3256 3756 3262 3762
rect 3314 3756 3320 3762
rect 7256 3756 7262 3762
rect 7314 3756 7320 3762
rect 11256 3756 11262 3762
rect 11314 3756 11320 3762
rect 15256 3756 15262 3762
rect 15314 3756 15320 3762
rect 19256 3756 19262 3762
rect 19314 3756 19320 3762
rect 23256 3756 23262 3762
rect 23314 3756 23320 3762
rect 27256 3756 27262 3762
rect 27314 3756 27320 3762
rect 31256 3756 31262 3762
rect 31314 3756 31320 3762
rect 35256 3756 35262 3762
rect 35314 3756 35320 3762
rect 39256 3756 39262 3762
rect 39314 3756 39320 3762
rect 3262 3750 3268 3756
rect 3308 3750 3314 3756
rect 7262 3750 7268 3756
rect 7308 3750 7314 3756
rect 11262 3750 11268 3756
rect 11308 3750 11314 3756
rect 15262 3750 15268 3756
rect 15308 3750 15314 3756
rect 19262 3750 19268 3756
rect 19308 3750 19314 3756
rect 23262 3750 23268 3756
rect 23308 3750 23314 3756
rect 27262 3750 27268 3756
rect 27308 3750 27314 3756
rect 31262 3750 31268 3756
rect 31308 3750 31314 3756
rect 35262 3750 35268 3756
rect 35308 3750 35314 3756
rect 39262 3750 39268 3756
rect 39308 3750 39314 3756
rect 2386 3296 2626 3320
rect 2386 3104 2410 3296
rect 2602 3104 2626 3296
rect 2386 3080 2626 3104
rect 6386 3296 6626 3320
rect 6386 3104 6410 3296
rect 6602 3104 6626 3296
rect 6386 3080 6626 3104
rect 10386 3296 10626 3320
rect 10386 3104 10410 3296
rect 10602 3104 10626 3296
rect 10386 3080 10626 3104
rect 14386 3296 14626 3320
rect 14386 3104 14410 3296
rect 14602 3104 14626 3296
rect 14386 3080 14626 3104
rect 18386 3296 18626 3320
rect 18386 3104 18410 3296
rect 18602 3104 18626 3296
rect 18386 3080 18626 3104
rect 22386 3296 22626 3320
rect 22386 3104 22410 3296
rect 22602 3104 22626 3296
rect 22386 3080 22626 3104
rect 26386 3296 26626 3320
rect 26386 3104 26410 3296
rect 26602 3104 26626 3296
rect 26386 3080 26626 3104
rect 30386 3296 30626 3320
rect 30386 3104 30410 3296
rect 30602 3104 30626 3296
rect 30386 3080 30626 3104
rect 34386 3296 34626 3320
rect 34386 3104 34410 3296
rect 34602 3104 34626 3296
rect 34386 3080 34626 3104
rect 38386 3296 38626 3320
rect 38386 3104 38410 3296
rect 38602 3104 38626 3296
rect 38386 3080 38626 3104
rect 1982 2160 2302 2230
rect 366 1916 606 1940
rect 366 1724 390 1916
rect 582 1724 606 1916
rect 1982 1920 2006 2160
rect 2232 1920 2246 2160
rect 2256 1920 2302 2160
rect 5982 2160 6302 2230
rect 1982 1896 2302 1920
rect 4366 1916 4606 1940
rect 366 1700 606 1724
rect 4366 1724 4390 1916
rect 4582 1724 4606 1916
rect 5982 1920 6006 2160
rect 6232 1920 6246 2160
rect 6256 1920 6302 2160
rect 9982 2160 10302 2230
rect 5982 1896 6302 1920
rect 8366 1916 8606 1940
rect 2852 1709 2996 1714
rect 2852 1639 2857 1709
rect 2991 1639 2996 1709
rect 4366 1700 4606 1724
rect 8366 1724 8390 1916
rect 8582 1724 8606 1916
rect 9982 1920 10006 2160
rect 10232 1920 10246 2160
rect 10256 1920 10302 2160
rect 13982 2160 14302 2230
rect 9982 1896 10302 1920
rect 12366 1916 12606 1940
rect 6852 1709 6996 1714
rect 2852 1634 2996 1639
rect 6852 1639 6857 1709
rect 6991 1639 6996 1709
rect 8366 1700 8606 1724
rect 12366 1724 12390 1916
rect 12582 1724 12606 1916
rect 13982 1920 14006 2160
rect 14232 1920 14246 2160
rect 14256 1920 14302 2160
rect 17982 2160 18302 2230
rect 13982 1896 14302 1920
rect 16366 1916 16606 1940
rect 10852 1709 10996 1714
rect 6852 1634 6996 1639
rect 10852 1639 10857 1709
rect 10991 1639 10996 1709
rect 12366 1700 12606 1724
rect 16366 1724 16390 1916
rect 16582 1724 16606 1916
rect 17982 1920 18006 2160
rect 18232 1920 18246 2160
rect 18256 1920 18302 2160
rect 21982 2160 22302 2230
rect 17982 1896 18302 1920
rect 20366 1916 20606 1940
rect 14852 1709 14996 1714
rect 10852 1634 10996 1639
rect 14852 1639 14857 1709
rect 14991 1639 14996 1709
rect 16366 1700 16606 1724
rect 20366 1724 20390 1916
rect 20582 1724 20606 1916
rect 21982 1920 22006 2160
rect 22232 1920 22246 2160
rect 22256 1920 22302 2160
rect 25982 2160 26302 2230
rect 21982 1896 22302 1920
rect 24366 1916 24606 1940
rect 18852 1709 18996 1714
rect 14852 1634 14996 1639
rect 18852 1639 18857 1709
rect 18991 1639 18996 1709
rect 20366 1700 20606 1724
rect 24366 1724 24390 1916
rect 24582 1724 24606 1916
rect 25982 1920 26006 2160
rect 26232 1920 26246 2160
rect 26256 1920 26302 2160
rect 29982 2160 30302 2230
rect 25982 1896 26302 1920
rect 28366 1916 28606 1940
rect 22852 1709 22996 1714
rect 18852 1634 18996 1639
rect 22852 1639 22857 1709
rect 22991 1639 22996 1709
rect 24366 1700 24606 1724
rect 28366 1724 28390 1916
rect 28582 1724 28606 1916
rect 29982 1920 30006 2160
rect 30232 1920 30246 2160
rect 30256 1920 30302 2160
rect 33982 2160 34302 2230
rect 29982 1896 30302 1920
rect 32366 1916 32606 1940
rect 26852 1709 26996 1714
rect 22852 1634 22996 1639
rect 26852 1639 26857 1709
rect 26991 1639 26996 1709
rect 28366 1700 28606 1724
rect 32366 1724 32390 1916
rect 32582 1724 32606 1916
rect 33982 1920 34006 2160
rect 34232 1920 34246 2160
rect 34256 1920 34302 2160
rect 37982 2160 38302 2230
rect 33982 1896 34302 1920
rect 36366 1916 36606 1940
rect 30852 1709 30996 1714
rect 26852 1634 26996 1639
rect 30852 1639 30857 1709
rect 30991 1639 30996 1709
rect 32366 1700 32606 1724
rect 36366 1724 36390 1916
rect 36582 1724 36606 1916
rect 37982 1920 38006 2160
rect 38232 1920 38246 2160
rect 38256 1920 38302 2160
rect 37982 1896 38302 1920
rect 34852 1709 34996 1714
rect 30852 1634 30996 1639
rect 34852 1639 34857 1709
rect 34991 1639 34996 1709
rect 36366 1700 36606 1724
rect 38852 1709 38996 1714
rect 34852 1634 34996 1639
rect 38852 1639 38857 1709
rect 38991 1639 38996 1709
rect 38852 1634 38996 1639
rect 2366 1559 2546 1560
rect 2366 1381 2367 1559
rect 2545 1381 2546 1559
rect 2366 1380 2546 1381
rect 6366 1559 6546 1560
rect 6366 1381 6367 1559
rect 6545 1381 6546 1559
rect 6366 1380 6546 1381
rect 10366 1559 10546 1560
rect 10366 1381 10367 1559
rect 10545 1381 10546 1559
rect 10366 1380 10546 1381
rect 14366 1559 14546 1560
rect 14366 1381 14367 1559
rect 14545 1381 14546 1559
rect 14366 1380 14546 1381
rect 18366 1559 18546 1560
rect 18366 1381 18367 1559
rect 18545 1381 18546 1559
rect 18366 1380 18546 1381
rect 22366 1559 22546 1560
rect 22366 1381 22367 1559
rect 22545 1381 22546 1559
rect 22366 1380 22546 1381
rect 26366 1559 26546 1560
rect 26366 1381 26367 1559
rect 26545 1381 26546 1559
rect 26366 1380 26546 1381
rect 30366 1559 30546 1560
rect 30366 1381 30367 1559
rect 30545 1381 30546 1559
rect 30366 1380 30546 1381
rect 34366 1559 34546 1560
rect 34366 1381 34367 1559
rect 34545 1381 34546 1559
rect 34366 1380 34546 1381
rect 38366 1559 38546 1560
rect 38366 1381 38367 1559
rect 38545 1381 38546 1559
rect 38366 1380 38546 1381
rect 366 1039 546 1040
rect 366 861 367 1039
rect 545 861 546 1039
rect 4366 1039 4546 1040
rect 3734 984 3740 990
rect 3780 984 3786 990
rect 3728 978 3734 984
rect 3786 978 3792 984
rect 3728 928 3734 934
rect 3786 928 3792 934
rect 3734 922 3740 928
rect 3780 922 3786 928
rect 366 860 546 861
rect 4366 861 4367 1039
rect 4545 861 4546 1039
rect 8366 1039 8546 1040
rect 7734 984 7740 990
rect 7780 984 7786 990
rect 7728 978 7734 984
rect 7786 978 7792 984
rect 7728 928 7734 934
rect 7786 928 7792 934
rect 7734 922 7740 928
rect 7780 922 7786 928
rect 4366 860 4546 861
rect 8366 861 8367 1039
rect 8545 861 8546 1039
rect 12366 1039 12546 1040
rect 11734 984 11740 990
rect 11780 984 11786 990
rect 11728 978 11734 984
rect 11786 978 11792 984
rect 11728 928 11734 934
rect 11786 928 11792 934
rect 11734 922 11740 928
rect 11780 922 11786 928
rect 8366 860 8546 861
rect 12366 861 12367 1039
rect 12545 861 12546 1039
rect 16366 1039 16546 1040
rect 15734 984 15740 990
rect 15780 984 15786 990
rect 15728 978 15734 984
rect 15786 978 15792 984
rect 15728 928 15734 934
rect 15786 928 15792 934
rect 15734 922 15740 928
rect 15780 922 15786 928
rect 12366 860 12546 861
rect 16366 861 16367 1039
rect 16545 861 16546 1039
rect 20366 1039 20546 1040
rect 19734 984 19740 990
rect 19780 984 19786 990
rect 19728 978 19734 984
rect 19786 978 19792 984
rect 19728 928 19734 934
rect 19786 928 19792 934
rect 19734 922 19740 928
rect 19780 922 19786 928
rect 16366 860 16546 861
rect 20366 861 20367 1039
rect 20545 861 20546 1039
rect 24366 1039 24546 1040
rect 23734 984 23740 990
rect 23780 984 23786 990
rect 23728 978 23734 984
rect 23786 978 23792 984
rect 23728 928 23734 934
rect 23786 928 23792 934
rect 23734 922 23740 928
rect 23780 922 23786 928
rect 20366 860 20546 861
rect 24366 861 24367 1039
rect 24545 861 24546 1039
rect 28366 1039 28546 1040
rect 27734 984 27740 990
rect 27780 984 27786 990
rect 27728 978 27734 984
rect 27786 978 27792 984
rect 27728 928 27734 934
rect 27786 928 27792 934
rect 27734 922 27740 928
rect 27780 922 27786 928
rect 24366 860 24546 861
rect 28366 861 28367 1039
rect 28545 861 28546 1039
rect 32366 1039 32546 1040
rect 31734 984 31740 990
rect 31780 984 31786 990
rect 31728 978 31734 984
rect 31786 978 31792 984
rect 31728 928 31734 934
rect 31786 928 31792 934
rect 31734 922 31740 928
rect 31780 922 31786 928
rect 28366 860 28546 861
rect 32366 861 32367 1039
rect 32545 861 32546 1039
rect 36366 1039 36546 1040
rect 35734 984 35740 990
rect 35780 984 35786 990
rect 35728 978 35734 984
rect 35786 978 35792 984
rect 35728 928 35734 934
rect 35786 928 35792 934
rect 35734 922 35740 928
rect 35780 922 35786 928
rect 32366 860 32546 861
rect 36366 861 36367 1039
rect 36545 861 36546 1039
rect 39734 984 39740 990
rect 39780 984 39786 990
rect 39728 978 39734 984
rect 39786 978 39792 984
rect 39728 928 39734 934
rect 39786 928 39792 934
rect 39734 922 39740 928
rect 39780 922 39786 928
rect 36366 860 36546 861
rect 3262 808 3268 814
rect 3308 808 3314 814
rect 7262 808 7268 814
rect 7308 808 7314 814
rect 11262 808 11268 814
rect 11308 808 11314 814
rect 15262 808 15268 814
rect 15308 808 15314 814
rect 19262 808 19268 814
rect 19308 808 19314 814
rect 23262 808 23268 814
rect 23308 808 23314 814
rect 27262 808 27268 814
rect 27308 808 27314 814
rect 31262 808 31268 814
rect 31308 808 31314 814
rect 35262 808 35268 814
rect 35308 808 35314 814
rect 39262 808 39268 814
rect 39308 808 39314 814
rect 3256 802 3262 808
rect 3314 802 3320 808
rect 7256 802 7262 808
rect 7314 802 7320 808
rect 11256 802 11262 808
rect 11314 802 11320 808
rect 15256 802 15262 808
rect 15314 802 15320 808
rect 19256 802 19262 808
rect 19314 802 19320 808
rect 23256 802 23262 808
rect 23314 802 23320 808
rect 27256 802 27262 808
rect 27314 802 27320 808
rect 31256 802 31262 808
rect 31314 802 31320 808
rect 35256 802 35262 808
rect 35314 802 35320 808
rect 39256 802 39262 808
rect 39314 802 39320 808
rect 3256 756 3262 762
rect 3314 756 3320 762
rect 7256 756 7262 762
rect 7314 756 7320 762
rect 11256 756 11262 762
rect 11314 756 11320 762
rect 15256 756 15262 762
rect 15314 756 15320 762
rect 19256 756 19262 762
rect 19314 756 19320 762
rect 23256 756 23262 762
rect 23314 756 23320 762
rect 27256 756 27262 762
rect 27314 756 27320 762
rect 31256 756 31262 762
rect 31314 756 31320 762
rect 35256 756 35262 762
rect 35314 756 35320 762
rect 39256 756 39262 762
rect 39314 756 39320 762
rect 3262 750 3268 756
rect 3308 750 3314 756
rect 7262 750 7268 756
rect 7308 750 7314 756
rect 11262 750 11268 756
rect 11308 750 11314 756
rect 15262 750 15268 756
rect 15308 750 15314 756
rect 19262 750 19268 756
rect 19308 750 19314 756
rect 23262 750 23268 756
rect 23308 750 23314 756
rect 27262 750 27268 756
rect 27308 750 27314 756
rect 31262 750 31268 756
rect 31308 750 31314 756
rect 35262 750 35268 756
rect 35308 750 35314 756
rect 39262 750 39268 756
rect 39308 750 39314 756
rect 2386 296 2626 320
rect 2386 104 2410 296
rect 2602 104 2626 296
rect 2386 80 2626 104
rect 6386 296 6626 320
rect 6386 104 6410 296
rect 6602 104 6626 296
rect 6386 80 6626 104
rect 10386 296 10626 320
rect 10386 104 10410 296
rect 10602 104 10626 296
rect 10386 80 10626 104
rect 14386 296 14626 320
rect 14386 104 14410 296
rect 14602 104 14626 296
rect 14386 80 14626 104
rect 18386 296 18626 320
rect 18386 104 18410 296
rect 18602 104 18626 296
rect 18386 80 18626 104
rect 22386 296 22626 320
rect 22386 104 22410 296
rect 22602 104 22626 296
rect 22386 80 22626 104
rect 26386 296 26626 320
rect 26386 104 26410 296
rect 26602 104 26626 296
rect 26386 80 26626 104
rect 30386 296 30626 320
rect 30386 104 30410 296
rect 30602 104 30626 296
rect 30386 80 30626 104
rect 34386 296 34626 320
rect 34386 104 34410 296
rect 34602 104 34626 296
rect 34386 80 34626 104
rect 38386 296 38626 320
rect 38386 104 38410 296
rect 38602 104 38626 296
rect 38386 80 38626 104
use fgcell_amp_nocap  fgcell_amp_nocap_0
array 0 9 4000 0 9 3000
timestamp 1717628967
transform 1 0 -140 0 1 7210
box 140 -7210 4106 -4964
<< end >>
