magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< error_p >>
rect 2240 28204 2480 28228
rect 2240 28142 2264 28204
rect 2456 28142 2480 28204
rect 2240 27988 2480 28142
rect 6240 28204 6480 28228
rect 6240 28142 6264 28204
rect 6456 28142 6480 28204
rect 6240 27988 6480 28142
rect 10240 28204 10480 28228
rect 10240 28142 10264 28204
rect 10456 28142 10480 28204
rect 10240 27988 10480 28142
rect 14240 28204 14480 28228
rect 14240 28142 14264 28204
rect 14456 28142 14480 28204
rect 14240 27988 14480 28142
rect 18240 28204 18480 28228
rect 18240 28142 18264 28204
rect 18456 28142 18480 28204
rect 18240 27988 18480 28142
rect 22240 28204 22480 28228
rect 22240 28142 22264 28204
rect 22456 28142 22480 28204
rect 22240 27988 22480 28142
rect 26240 28204 26480 28228
rect 26240 28142 26264 28204
rect 26456 28142 26480 28204
rect 26240 27988 26480 28142
rect 30240 28204 30480 28228
rect 30240 28142 30264 28204
rect 30456 28142 30480 28204
rect 30240 27988 30480 28142
rect 34240 28204 34480 28228
rect 34240 28142 34264 28204
rect 34456 28142 34480 28204
rect 34240 27988 34480 28142
rect 38240 28204 38480 28228
rect 38240 28142 38264 28204
rect 38456 28142 38480 28204
rect 38240 27988 38480 28142
rect 1934 27768 2254 27822
rect 360 27524 600 27548
rect 360 27332 384 27524
rect 576 27332 600 27524
rect 1934 27528 1960 27768
rect 2182 27528 2200 27768
rect 2206 27528 2254 27768
rect 3602 27771 3690 27776
rect 3602 27693 3607 27771
rect 3685 27693 3690 27771
rect 3602 27688 3690 27693
rect 5934 27768 6254 27822
rect 1934 27502 2254 27528
rect 4360 27524 4600 27548
rect 360 27308 600 27332
rect 4360 27332 4384 27524
rect 4576 27332 4600 27524
rect 5934 27528 5960 27768
rect 6182 27528 6200 27768
rect 6206 27528 6254 27768
rect 7602 27771 7690 27776
rect 7602 27693 7607 27771
rect 7685 27693 7690 27771
rect 7602 27688 7690 27693
rect 9934 27768 10254 27822
rect 5934 27502 6254 27528
rect 8360 27524 8600 27548
rect 2810 27319 2946 27324
rect 2810 27245 2815 27319
rect 2941 27245 2946 27319
rect 4360 27308 4600 27332
rect 8360 27332 8384 27524
rect 8576 27332 8600 27524
rect 9934 27528 9960 27768
rect 10182 27528 10200 27768
rect 10206 27528 10254 27768
rect 11602 27771 11690 27776
rect 11602 27693 11607 27771
rect 11685 27693 11690 27771
rect 11602 27688 11690 27693
rect 13934 27768 14254 27822
rect 9934 27502 10254 27528
rect 12360 27524 12600 27548
rect 6810 27319 6946 27324
rect 2810 27240 2946 27245
rect 6810 27245 6815 27319
rect 6941 27245 6946 27319
rect 8360 27308 8600 27332
rect 12360 27332 12384 27524
rect 12576 27332 12600 27524
rect 13934 27528 13960 27768
rect 14182 27528 14200 27768
rect 14206 27528 14254 27768
rect 15602 27771 15690 27776
rect 15602 27693 15607 27771
rect 15685 27693 15690 27771
rect 15602 27688 15690 27693
rect 17934 27768 18254 27822
rect 13934 27502 14254 27528
rect 16360 27524 16600 27548
rect 10810 27319 10946 27324
rect 6810 27240 6946 27245
rect 10810 27245 10815 27319
rect 10941 27245 10946 27319
rect 12360 27308 12600 27332
rect 16360 27332 16384 27524
rect 16576 27332 16600 27524
rect 17934 27528 17960 27768
rect 18182 27528 18200 27768
rect 18206 27528 18254 27768
rect 19602 27771 19690 27776
rect 19602 27693 19607 27771
rect 19685 27693 19690 27771
rect 19602 27688 19690 27693
rect 21934 27768 22254 27822
rect 17934 27502 18254 27528
rect 20360 27524 20600 27548
rect 14810 27319 14946 27324
rect 10810 27240 10946 27245
rect 14810 27245 14815 27319
rect 14941 27245 14946 27319
rect 16360 27308 16600 27332
rect 20360 27332 20384 27524
rect 20576 27332 20600 27524
rect 21934 27528 21960 27768
rect 22182 27528 22200 27768
rect 22206 27528 22254 27768
rect 23602 27771 23690 27776
rect 23602 27693 23607 27771
rect 23685 27693 23690 27771
rect 23602 27688 23690 27693
rect 25934 27768 26254 27822
rect 21934 27502 22254 27528
rect 24360 27524 24600 27548
rect 18810 27319 18946 27324
rect 14810 27240 14946 27245
rect 18810 27245 18815 27319
rect 18941 27245 18946 27319
rect 20360 27308 20600 27332
rect 24360 27332 24384 27524
rect 24576 27332 24600 27524
rect 25934 27528 25960 27768
rect 26182 27528 26200 27768
rect 26206 27528 26254 27768
rect 27602 27771 27690 27776
rect 27602 27693 27607 27771
rect 27685 27693 27690 27771
rect 27602 27688 27690 27693
rect 29934 27768 30254 27822
rect 25934 27502 26254 27528
rect 28360 27524 28600 27548
rect 22810 27319 22946 27324
rect 18810 27240 18946 27245
rect 22810 27245 22815 27319
rect 22941 27245 22946 27319
rect 24360 27308 24600 27332
rect 28360 27332 28384 27524
rect 28576 27332 28600 27524
rect 29934 27528 29960 27768
rect 30182 27528 30200 27768
rect 30206 27528 30254 27768
rect 31602 27771 31690 27776
rect 31602 27693 31607 27771
rect 31685 27693 31690 27771
rect 31602 27688 31690 27693
rect 33934 27768 34254 27822
rect 29934 27502 30254 27528
rect 32360 27524 32600 27548
rect 26810 27319 26946 27324
rect 22810 27240 22946 27245
rect 26810 27245 26815 27319
rect 26941 27245 26946 27319
rect 28360 27308 28600 27332
rect 32360 27332 32384 27524
rect 32576 27332 32600 27524
rect 33934 27528 33960 27768
rect 34182 27528 34200 27768
rect 34206 27528 34254 27768
rect 35602 27771 35690 27776
rect 35602 27693 35607 27771
rect 35685 27693 35690 27771
rect 35602 27688 35690 27693
rect 37934 27768 38254 27822
rect 33934 27502 34254 27528
rect 36360 27524 36600 27548
rect 30810 27319 30946 27324
rect 26810 27240 26946 27245
rect 30810 27245 30815 27319
rect 30941 27245 30946 27319
rect 32360 27308 32600 27332
rect 36360 27332 36384 27524
rect 36576 27332 36600 27524
rect 37934 27528 37960 27768
rect 38182 27528 38200 27768
rect 38206 27528 38254 27768
rect 39602 27771 39690 27776
rect 39602 27693 39607 27771
rect 39685 27693 39690 27771
rect 39602 27688 39690 27693
rect 37934 27502 38254 27528
rect 34810 27319 34946 27324
rect 30810 27240 30946 27245
rect 34810 27245 34815 27319
rect 34941 27245 34946 27319
rect 36360 27308 36600 27332
rect 38810 27319 38946 27324
rect 34810 27240 34946 27245
rect 38810 27245 38815 27319
rect 38941 27245 38946 27319
rect 38810 27240 38946 27245
rect 2338 27181 2518 27182
rect 2338 27003 2339 27181
rect 2517 27003 2518 27181
rect 2338 27002 2518 27003
rect 6338 27181 6518 27182
rect 6338 27003 6339 27181
rect 6517 27003 6518 27181
rect 6338 27002 6518 27003
rect 10338 27181 10518 27182
rect 10338 27003 10339 27181
rect 10517 27003 10518 27181
rect 10338 27002 10518 27003
rect 14338 27181 14518 27182
rect 14338 27003 14339 27181
rect 14517 27003 14518 27181
rect 14338 27002 14518 27003
rect 18338 27181 18518 27182
rect 18338 27003 18339 27181
rect 18517 27003 18518 27181
rect 18338 27002 18518 27003
rect 22338 27181 22518 27182
rect 22338 27003 22339 27181
rect 22517 27003 22518 27181
rect 22338 27002 22518 27003
rect 26338 27181 26518 27182
rect 26338 27003 26339 27181
rect 26517 27003 26518 27181
rect 26338 27002 26518 27003
rect 30338 27181 30518 27182
rect 30338 27003 30339 27181
rect 30517 27003 30518 27181
rect 30338 27002 30518 27003
rect 34338 27181 34518 27182
rect 34338 27003 34339 27181
rect 34517 27003 34518 27181
rect 34338 27002 34518 27003
rect 38338 27181 38518 27182
rect 38338 27003 38339 27181
rect 38517 27003 38518 27181
rect 38338 27002 38518 27003
rect 390 26607 570 26608
rect 390 26429 391 26607
rect 569 26429 570 26607
rect 3734 26604 3740 26610
rect 3780 26604 3786 26610
rect 4390 26607 4570 26608
rect 3728 26598 3734 26604
rect 3786 26598 3792 26604
rect 3728 26552 3734 26558
rect 3786 26552 3792 26558
rect 3734 26546 3740 26552
rect 3780 26546 3786 26552
rect 390 26428 570 26429
rect 4390 26429 4391 26607
rect 4569 26429 4570 26607
rect 7734 26604 7740 26610
rect 7780 26604 7786 26610
rect 8390 26607 8570 26608
rect 7728 26598 7734 26604
rect 7786 26598 7792 26604
rect 7728 26552 7734 26558
rect 7786 26552 7792 26558
rect 7734 26546 7740 26552
rect 7780 26546 7786 26552
rect 4390 26428 4570 26429
rect 8390 26429 8391 26607
rect 8569 26429 8570 26607
rect 11734 26604 11740 26610
rect 11780 26604 11786 26610
rect 12390 26607 12570 26608
rect 11728 26598 11734 26604
rect 11786 26598 11792 26604
rect 11728 26552 11734 26558
rect 11786 26552 11792 26558
rect 11734 26546 11740 26552
rect 11780 26546 11786 26552
rect 8390 26428 8570 26429
rect 12390 26429 12391 26607
rect 12569 26429 12570 26607
rect 15734 26604 15740 26610
rect 15780 26604 15786 26610
rect 16390 26607 16570 26608
rect 15728 26598 15734 26604
rect 15786 26598 15792 26604
rect 15728 26552 15734 26558
rect 15786 26552 15792 26558
rect 15734 26546 15740 26552
rect 15780 26546 15786 26552
rect 12390 26428 12570 26429
rect 16390 26429 16391 26607
rect 16569 26429 16570 26607
rect 19734 26604 19740 26610
rect 19780 26604 19786 26610
rect 20390 26607 20570 26608
rect 19728 26598 19734 26604
rect 19786 26598 19792 26604
rect 19728 26552 19734 26558
rect 19786 26552 19792 26558
rect 19734 26546 19740 26552
rect 19780 26546 19786 26552
rect 16390 26428 16570 26429
rect 20390 26429 20391 26607
rect 20569 26429 20570 26607
rect 23734 26604 23740 26610
rect 23780 26604 23786 26610
rect 24390 26607 24570 26608
rect 23728 26598 23734 26604
rect 23786 26598 23792 26604
rect 23728 26552 23734 26558
rect 23786 26552 23792 26558
rect 23734 26546 23740 26552
rect 23780 26546 23786 26552
rect 20390 26428 20570 26429
rect 24390 26429 24391 26607
rect 24569 26429 24570 26607
rect 27734 26604 27740 26610
rect 27780 26604 27786 26610
rect 28390 26607 28570 26608
rect 27728 26598 27734 26604
rect 27786 26598 27792 26604
rect 27728 26552 27734 26558
rect 27786 26552 27792 26558
rect 27734 26546 27740 26552
rect 27780 26546 27786 26552
rect 24390 26428 24570 26429
rect 28390 26429 28391 26607
rect 28569 26429 28570 26607
rect 31734 26604 31740 26610
rect 31780 26604 31786 26610
rect 32390 26607 32570 26608
rect 31728 26598 31734 26604
rect 31786 26598 31792 26604
rect 31728 26552 31734 26558
rect 31786 26552 31792 26558
rect 31734 26546 31740 26552
rect 31780 26546 31786 26552
rect 28390 26428 28570 26429
rect 32390 26429 32391 26607
rect 32569 26429 32570 26607
rect 35734 26604 35740 26610
rect 35780 26604 35786 26610
rect 36390 26607 36570 26608
rect 35728 26598 35734 26604
rect 35786 26598 35792 26604
rect 35728 26552 35734 26558
rect 35786 26552 35792 26558
rect 35734 26546 35740 26552
rect 35780 26546 35786 26552
rect 32390 26428 32570 26429
rect 36390 26429 36391 26607
rect 36569 26429 36570 26607
rect 39734 26604 39740 26610
rect 39780 26604 39786 26610
rect 39728 26598 39734 26604
rect 39786 26598 39792 26604
rect 39728 26552 39734 26558
rect 39786 26552 39792 26558
rect 39734 26546 39740 26552
rect 39780 26546 39786 26552
rect 36390 26428 36570 26429
rect 3262 26416 3268 26422
rect 3308 26416 3314 26422
rect 7262 26416 7268 26422
rect 7308 26416 7314 26422
rect 11262 26416 11268 26422
rect 11308 26416 11314 26422
rect 15262 26416 15268 26422
rect 15308 26416 15314 26422
rect 19262 26416 19268 26422
rect 19308 26416 19314 26422
rect 23262 26416 23268 26422
rect 23308 26416 23314 26422
rect 27262 26416 27268 26422
rect 27308 26416 27314 26422
rect 31262 26416 31268 26422
rect 31308 26416 31314 26422
rect 35262 26416 35268 26422
rect 35308 26416 35314 26422
rect 39262 26416 39268 26422
rect 39308 26416 39314 26422
rect 3256 26410 3262 26416
rect 3314 26410 3320 26416
rect 7256 26410 7262 26416
rect 7314 26410 7320 26416
rect 11256 26410 11262 26416
rect 11314 26410 11320 26416
rect 15256 26410 15262 26416
rect 15314 26410 15320 26416
rect 19256 26410 19262 26416
rect 19314 26410 19320 26416
rect 23256 26410 23262 26416
rect 23314 26410 23320 26416
rect 27256 26410 27262 26416
rect 27314 26410 27320 26416
rect 31256 26410 31262 26416
rect 31314 26410 31320 26416
rect 35256 26410 35262 26416
rect 35314 26410 35320 26416
rect 39256 26410 39262 26416
rect 39314 26410 39320 26416
rect 3256 26364 3262 26370
rect 3314 26364 3320 26370
rect 7256 26364 7262 26370
rect 7314 26364 7320 26370
rect 11256 26364 11262 26370
rect 11314 26364 11320 26370
rect 15256 26364 15262 26370
rect 15314 26364 15320 26370
rect 19256 26364 19262 26370
rect 19314 26364 19320 26370
rect 23256 26364 23262 26370
rect 23314 26364 23320 26370
rect 27256 26364 27262 26370
rect 27314 26364 27320 26370
rect 31256 26364 31262 26370
rect 31314 26364 31320 26370
rect 35256 26364 35262 26370
rect 35314 26364 35320 26370
rect 39256 26364 39262 26370
rect 39314 26364 39320 26370
rect 3262 26358 3268 26364
rect 3308 26358 3314 26364
rect 7262 26358 7268 26364
rect 7308 26358 7314 26364
rect 11262 26358 11268 26364
rect 11308 26358 11314 26364
rect 15262 26358 15268 26364
rect 15308 26358 15314 26364
rect 19262 26358 19268 26364
rect 19308 26358 19314 26364
rect 23262 26358 23268 26364
rect 23308 26358 23314 26364
rect 27262 26358 27268 26364
rect 27308 26358 27314 26364
rect 31262 26358 31268 26364
rect 31308 26358 31314 26364
rect 35262 26358 35268 26364
rect 35308 26358 35314 26364
rect 39262 26358 39268 26364
rect 39308 26358 39314 26364
rect 2240 25904 2480 25928
rect 2240 25712 2264 25904
rect 2456 25712 2480 25904
rect 2240 25688 2480 25712
rect 6240 25904 6480 25928
rect 6240 25712 6264 25904
rect 6456 25712 6480 25904
rect 6240 25688 6480 25712
rect 10240 25904 10480 25928
rect 10240 25712 10264 25904
rect 10456 25712 10480 25904
rect 10240 25688 10480 25712
rect 14240 25904 14480 25928
rect 14240 25712 14264 25904
rect 14456 25712 14480 25904
rect 14240 25688 14480 25712
rect 18240 25904 18480 25928
rect 18240 25712 18264 25904
rect 18456 25712 18480 25904
rect 18240 25688 18480 25712
rect 22240 25904 22480 25928
rect 22240 25712 22264 25904
rect 22456 25712 22480 25904
rect 22240 25688 22480 25712
rect 26240 25904 26480 25928
rect 26240 25712 26264 25904
rect 26456 25712 26480 25904
rect 26240 25688 26480 25712
rect 30240 25904 30480 25928
rect 30240 25712 30264 25904
rect 30456 25712 30480 25904
rect 30240 25688 30480 25712
rect 34240 25904 34480 25928
rect 34240 25712 34264 25904
rect 34456 25712 34480 25904
rect 34240 25688 34480 25712
rect 38240 25904 38480 25928
rect 38240 25712 38264 25904
rect 38456 25712 38480 25904
rect 38240 25688 38480 25712
rect 2240 25204 2480 25228
rect 2240 25142 2264 25204
rect 2456 25142 2480 25204
rect 2240 24988 2480 25142
rect 6240 25204 6480 25228
rect 6240 25142 6264 25204
rect 6456 25142 6480 25204
rect 6240 24988 6480 25142
rect 10240 25204 10480 25228
rect 10240 25142 10264 25204
rect 10456 25142 10480 25204
rect 10240 24988 10480 25142
rect 14240 25204 14480 25228
rect 14240 25142 14264 25204
rect 14456 25142 14480 25204
rect 14240 24988 14480 25142
rect 18240 25204 18480 25228
rect 18240 25142 18264 25204
rect 18456 25142 18480 25204
rect 18240 24988 18480 25142
rect 22240 25204 22480 25228
rect 22240 25142 22264 25204
rect 22456 25142 22480 25204
rect 22240 24988 22480 25142
rect 26240 25204 26480 25228
rect 26240 25142 26264 25204
rect 26456 25142 26480 25204
rect 26240 24988 26480 25142
rect 30240 25204 30480 25228
rect 30240 25142 30264 25204
rect 30456 25142 30480 25204
rect 30240 24988 30480 25142
rect 34240 25204 34480 25228
rect 34240 25142 34264 25204
rect 34456 25142 34480 25204
rect 34240 24988 34480 25142
rect 38240 25204 38480 25228
rect 38240 25142 38264 25204
rect 38456 25142 38480 25204
rect 38240 24988 38480 25142
rect 1934 24768 2254 24822
rect 360 24524 600 24548
rect 360 24332 384 24524
rect 576 24332 600 24524
rect 1934 24528 1960 24768
rect 2182 24528 2200 24768
rect 2206 24528 2254 24768
rect 3602 24771 3690 24776
rect 3602 24693 3607 24771
rect 3685 24693 3690 24771
rect 3602 24688 3690 24693
rect 5934 24768 6254 24822
rect 1934 24502 2254 24528
rect 4360 24524 4600 24548
rect 360 24308 600 24332
rect 4360 24332 4384 24524
rect 4576 24332 4600 24524
rect 5934 24528 5960 24768
rect 6182 24528 6200 24768
rect 6206 24528 6254 24768
rect 7602 24771 7690 24776
rect 7602 24693 7607 24771
rect 7685 24693 7690 24771
rect 7602 24688 7690 24693
rect 9934 24768 10254 24822
rect 5934 24502 6254 24528
rect 8360 24524 8600 24548
rect 2810 24319 2946 24324
rect 2810 24245 2815 24319
rect 2941 24245 2946 24319
rect 4360 24308 4600 24332
rect 8360 24332 8384 24524
rect 8576 24332 8600 24524
rect 9934 24528 9960 24768
rect 10182 24528 10200 24768
rect 10206 24528 10254 24768
rect 11602 24771 11690 24776
rect 11602 24693 11607 24771
rect 11685 24693 11690 24771
rect 11602 24688 11690 24693
rect 13934 24768 14254 24822
rect 9934 24502 10254 24528
rect 12360 24524 12600 24548
rect 6810 24319 6946 24324
rect 2810 24240 2946 24245
rect 6810 24245 6815 24319
rect 6941 24245 6946 24319
rect 8360 24308 8600 24332
rect 12360 24332 12384 24524
rect 12576 24332 12600 24524
rect 13934 24528 13960 24768
rect 14182 24528 14200 24768
rect 14206 24528 14254 24768
rect 15602 24771 15690 24776
rect 15602 24693 15607 24771
rect 15685 24693 15690 24771
rect 15602 24688 15690 24693
rect 17934 24768 18254 24822
rect 13934 24502 14254 24528
rect 16360 24524 16600 24548
rect 10810 24319 10946 24324
rect 6810 24240 6946 24245
rect 10810 24245 10815 24319
rect 10941 24245 10946 24319
rect 12360 24308 12600 24332
rect 16360 24332 16384 24524
rect 16576 24332 16600 24524
rect 17934 24528 17960 24768
rect 18182 24528 18200 24768
rect 18206 24528 18254 24768
rect 19602 24771 19690 24776
rect 19602 24693 19607 24771
rect 19685 24693 19690 24771
rect 19602 24688 19690 24693
rect 21934 24768 22254 24822
rect 17934 24502 18254 24528
rect 20360 24524 20600 24548
rect 14810 24319 14946 24324
rect 10810 24240 10946 24245
rect 14810 24245 14815 24319
rect 14941 24245 14946 24319
rect 16360 24308 16600 24332
rect 20360 24332 20384 24524
rect 20576 24332 20600 24524
rect 21934 24528 21960 24768
rect 22182 24528 22200 24768
rect 22206 24528 22254 24768
rect 23602 24771 23690 24776
rect 23602 24693 23607 24771
rect 23685 24693 23690 24771
rect 23602 24688 23690 24693
rect 25934 24768 26254 24822
rect 21934 24502 22254 24528
rect 24360 24524 24600 24548
rect 18810 24319 18946 24324
rect 14810 24240 14946 24245
rect 18810 24245 18815 24319
rect 18941 24245 18946 24319
rect 20360 24308 20600 24332
rect 24360 24332 24384 24524
rect 24576 24332 24600 24524
rect 25934 24528 25960 24768
rect 26182 24528 26200 24768
rect 26206 24528 26254 24768
rect 27602 24771 27690 24776
rect 27602 24693 27607 24771
rect 27685 24693 27690 24771
rect 27602 24688 27690 24693
rect 29934 24768 30254 24822
rect 25934 24502 26254 24528
rect 28360 24524 28600 24548
rect 22810 24319 22946 24324
rect 18810 24240 18946 24245
rect 22810 24245 22815 24319
rect 22941 24245 22946 24319
rect 24360 24308 24600 24332
rect 28360 24332 28384 24524
rect 28576 24332 28600 24524
rect 29934 24528 29960 24768
rect 30182 24528 30200 24768
rect 30206 24528 30254 24768
rect 31602 24771 31690 24776
rect 31602 24693 31607 24771
rect 31685 24693 31690 24771
rect 31602 24688 31690 24693
rect 33934 24768 34254 24822
rect 29934 24502 30254 24528
rect 32360 24524 32600 24548
rect 26810 24319 26946 24324
rect 22810 24240 22946 24245
rect 26810 24245 26815 24319
rect 26941 24245 26946 24319
rect 28360 24308 28600 24332
rect 32360 24332 32384 24524
rect 32576 24332 32600 24524
rect 33934 24528 33960 24768
rect 34182 24528 34200 24768
rect 34206 24528 34254 24768
rect 35602 24771 35690 24776
rect 35602 24693 35607 24771
rect 35685 24693 35690 24771
rect 35602 24688 35690 24693
rect 37934 24768 38254 24822
rect 33934 24502 34254 24528
rect 36360 24524 36600 24548
rect 30810 24319 30946 24324
rect 26810 24240 26946 24245
rect 30810 24245 30815 24319
rect 30941 24245 30946 24319
rect 32360 24308 32600 24332
rect 36360 24332 36384 24524
rect 36576 24332 36600 24524
rect 37934 24528 37960 24768
rect 38182 24528 38200 24768
rect 38206 24528 38254 24768
rect 39602 24771 39690 24776
rect 39602 24693 39607 24771
rect 39685 24693 39690 24771
rect 39602 24688 39690 24693
rect 37934 24502 38254 24528
rect 34810 24319 34946 24324
rect 30810 24240 30946 24245
rect 34810 24245 34815 24319
rect 34941 24245 34946 24319
rect 36360 24308 36600 24332
rect 38810 24319 38946 24324
rect 34810 24240 34946 24245
rect 38810 24245 38815 24319
rect 38941 24245 38946 24319
rect 38810 24240 38946 24245
rect 2338 24181 2518 24182
rect 2338 24003 2339 24181
rect 2517 24003 2518 24181
rect 2338 24002 2518 24003
rect 6338 24181 6518 24182
rect 6338 24003 6339 24181
rect 6517 24003 6518 24181
rect 6338 24002 6518 24003
rect 10338 24181 10518 24182
rect 10338 24003 10339 24181
rect 10517 24003 10518 24181
rect 10338 24002 10518 24003
rect 14338 24181 14518 24182
rect 14338 24003 14339 24181
rect 14517 24003 14518 24181
rect 14338 24002 14518 24003
rect 18338 24181 18518 24182
rect 18338 24003 18339 24181
rect 18517 24003 18518 24181
rect 18338 24002 18518 24003
rect 22338 24181 22518 24182
rect 22338 24003 22339 24181
rect 22517 24003 22518 24181
rect 22338 24002 22518 24003
rect 26338 24181 26518 24182
rect 26338 24003 26339 24181
rect 26517 24003 26518 24181
rect 26338 24002 26518 24003
rect 30338 24181 30518 24182
rect 30338 24003 30339 24181
rect 30517 24003 30518 24181
rect 30338 24002 30518 24003
rect 34338 24181 34518 24182
rect 34338 24003 34339 24181
rect 34517 24003 34518 24181
rect 34338 24002 34518 24003
rect 38338 24181 38518 24182
rect 38338 24003 38339 24181
rect 38517 24003 38518 24181
rect 38338 24002 38518 24003
rect 390 23607 570 23608
rect 390 23429 391 23607
rect 569 23429 570 23607
rect 3734 23604 3740 23610
rect 3780 23604 3786 23610
rect 4390 23607 4570 23608
rect 3728 23598 3734 23604
rect 3786 23598 3792 23604
rect 3728 23552 3734 23558
rect 3786 23552 3792 23558
rect 3734 23546 3740 23552
rect 3780 23546 3786 23552
rect 390 23428 570 23429
rect 4390 23429 4391 23607
rect 4569 23429 4570 23607
rect 7734 23604 7740 23610
rect 7780 23604 7786 23610
rect 8390 23607 8570 23608
rect 7728 23598 7734 23604
rect 7786 23598 7792 23604
rect 7728 23552 7734 23558
rect 7786 23552 7792 23558
rect 7734 23546 7740 23552
rect 7780 23546 7786 23552
rect 4390 23428 4570 23429
rect 8390 23429 8391 23607
rect 8569 23429 8570 23607
rect 11734 23604 11740 23610
rect 11780 23604 11786 23610
rect 12390 23607 12570 23608
rect 11728 23598 11734 23604
rect 11786 23598 11792 23604
rect 11728 23552 11734 23558
rect 11786 23552 11792 23558
rect 11734 23546 11740 23552
rect 11780 23546 11786 23552
rect 8390 23428 8570 23429
rect 12390 23429 12391 23607
rect 12569 23429 12570 23607
rect 15734 23604 15740 23610
rect 15780 23604 15786 23610
rect 16390 23607 16570 23608
rect 15728 23598 15734 23604
rect 15786 23598 15792 23604
rect 15728 23552 15734 23558
rect 15786 23552 15792 23558
rect 15734 23546 15740 23552
rect 15780 23546 15786 23552
rect 12390 23428 12570 23429
rect 16390 23429 16391 23607
rect 16569 23429 16570 23607
rect 19734 23604 19740 23610
rect 19780 23604 19786 23610
rect 20390 23607 20570 23608
rect 19728 23598 19734 23604
rect 19786 23598 19792 23604
rect 19728 23552 19734 23558
rect 19786 23552 19792 23558
rect 19734 23546 19740 23552
rect 19780 23546 19786 23552
rect 16390 23428 16570 23429
rect 20390 23429 20391 23607
rect 20569 23429 20570 23607
rect 23734 23604 23740 23610
rect 23780 23604 23786 23610
rect 24390 23607 24570 23608
rect 23728 23598 23734 23604
rect 23786 23598 23792 23604
rect 23728 23552 23734 23558
rect 23786 23552 23792 23558
rect 23734 23546 23740 23552
rect 23780 23546 23786 23552
rect 20390 23428 20570 23429
rect 24390 23429 24391 23607
rect 24569 23429 24570 23607
rect 27734 23604 27740 23610
rect 27780 23604 27786 23610
rect 28390 23607 28570 23608
rect 27728 23598 27734 23604
rect 27786 23598 27792 23604
rect 27728 23552 27734 23558
rect 27786 23552 27792 23558
rect 27734 23546 27740 23552
rect 27780 23546 27786 23552
rect 24390 23428 24570 23429
rect 28390 23429 28391 23607
rect 28569 23429 28570 23607
rect 31734 23604 31740 23610
rect 31780 23604 31786 23610
rect 32390 23607 32570 23608
rect 31728 23598 31734 23604
rect 31786 23598 31792 23604
rect 31728 23552 31734 23558
rect 31786 23552 31792 23558
rect 31734 23546 31740 23552
rect 31780 23546 31786 23552
rect 28390 23428 28570 23429
rect 32390 23429 32391 23607
rect 32569 23429 32570 23607
rect 35734 23604 35740 23610
rect 35780 23604 35786 23610
rect 36390 23607 36570 23608
rect 35728 23598 35734 23604
rect 35786 23598 35792 23604
rect 35728 23552 35734 23558
rect 35786 23552 35792 23558
rect 35734 23546 35740 23552
rect 35780 23546 35786 23552
rect 32390 23428 32570 23429
rect 36390 23429 36391 23607
rect 36569 23429 36570 23607
rect 39734 23604 39740 23610
rect 39780 23604 39786 23610
rect 39728 23598 39734 23604
rect 39786 23598 39792 23604
rect 39728 23552 39734 23558
rect 39786 23552 39792 23558
rect 39734 23546 39740 23552
rect 39780 23546 39786 23552
rect 36390 23428 36570 23429
rect 3262 23416 3268 23422
rect 3308 23416 3314 23422
rect 7262 23416 7268 23422
rect 7308 23416 7314 23422
rect 11262 23416 11268 23422
rect 11308 23416 11314 23422
rect 15262 23416 15268 23422
rect 15308 23416 15314 23422
rect 19262 23416 19268 23422
rect 19308 23416 19314 23422
rect 23262 23416 23268 23422
rect 23308 23416 23314 23422
rect 27262 23416 27268 23422
rect 27308 23416 27314 23422
rect 31262 23416 31268 23422
rect 31308 23416 31314 23422
rect 35262 23416 35268 23422
rect 35308 23416 35314 23422
rect 39262 23416 39268 23422
rect 39308 23416 39314 23422
rect 3256 23410 3262 23416
rect 3314 23410 3320 23416
rect 7256 23410 7262 23416
rect 7314 23410 7320 23416
rect 11256 23410 11262 23416
rect 11314 23410 11320 23416
rect 15256 23410 15262 23416
rect 15314 23410 15320 23416
rect 19256 23410 19262 23416
rect 19314 23410 19320 23416
rect 23256 23410 23262 23416
rect 23314 23410 23320 23416
rect 27256 23410 27262 23416
rect 27314 23410 27320 23416
rect 31256 23410 31262 23416
rect 31314 23410 31320 23416
rect 35256 23410 35262 23416
rect 35314 23410 35320 23416
rect 39256 23410 39262 23416
rect 39314 23410 39320 23416
rect 3256 23364 3262 23370
rect 3314 23364 3320 23370
rect 7256 23364 7262 23370
rect 7314 23364 7320 23370
rect 11256 23364 11262 23370
rect 11314 23364 11320 23370
rect 15256 23364 15262 23370
rect 15314 23364 15320 23370
rect 19256 23364 19262 23370
rect 19314 23364 19320 23370
rect 23256 23364 23262 23370
rect 23314 23364 23320 23370
rect 27256 23364 27262 23370
rect 27314 23364 27320 23370
rect 31256 23364 31262 23370
rect 31314 23364 31320 23370
rect 35256 23364 35262 23370
rect 35314 23364 35320 23370
rect 39256 23364 39262 23370
rect 39314 23364 39320 23370
rect 3262 23358 3268 23364
rect 3308 23358 3314 23364
rect 7262 23358 7268 23364
rect 7308 23358 7314 23364
rect 11262 23358 11268 23364
rect 11308 23358 11314 23364
rect 15262 23358 15268 23364
rect 15308 23358 15314 23364
rect 19262 23358 19268 23364
rect 19308 23358 19314 23364
rect 23262 23358 23268 23364
rect 23308 23358 23314 23364
rect 27262 23358 27268 23364
rect 27308 23358 27314 23364
rect 31262 23358 31268 23364
rect 31308 23358 31314 23364
rect 35262 23358 35268 23364
rect 35308 23358 35314 23364
rect 39262 23358 39268 23364
rect 39308 23358 39314 23364
rect 2240 22904 2480 22928
rect 2240 22712 2264 22904
rect 2456 22712 2480 22904
rect 2240 22688 2480 22712
rect 6240 22904 6480 22928
rect 6240 22712 6264 22904
rect 6456 22712 6480 22904
rect 6240 22688 6480 22712
rect 10240 22904 10480 22928
rect 10240 22712 10264 22904
rect 10456 22712 10480 22904
rect 10240 22688 10480 22712
rect 14240 22904 14480 22928
rect 14240 22712 14264 22904
rect 14456 22712 14480 22904
rect 14240 22688 14480 22712
rect 18240 22904 18480 22928
rect 18240 22712 18264 22904
rect 18456 22712 18480 22904
rect 18240 22688 18480 22712
rect 22240 22904 22480 22928
rect 22240 22712 22264 22904
rect 22456 22712 22480 22904
rect 22240 22688 22480 22712
rect 26240 22904 26480 22928
rect 26240 22712 26264 22904
rect 26456 22712 26480 22904
rect 26240 22688 26480 22712
rect 30240 22904 30480 22928
rect 30240 22712 30264 22904
rect 30456 22712 30480 22904
rect 30240 22688 30480 22712
rect 34240 22904 34480 22928
rect 34240 22712 34264 22904
rect 34456 22712 34480 22904
rect 34240 22688 34480 22712
rect 38240 22904 38480 22928
rect 38240 22712 38264 22904
rect 38456 22712 38480 22904
rect 38240 22688 38480 22712
rect 2240 22204 2480 22228
rect 2240 22142 2264 22204
rect 2456 22142 2480 22204
rect 2240 21988 2480 22142
rect 6240 22204 6480 22228
rect 6240 22142 6264 22204
rect 6456 22142 6480 22204
rect 6240 21988 6480 22142
rect 10240 22204 10480 22228
rect 10240 22142 10264 22204
rect 10456 22142 10480 22204
rect 10240 21988 10480 22142
rect 14240 22204 14480 22228
rect 14240 22142 14264 22204
rect 14456 22142 14480 22204
rect 14240 21988 14480 22142
rect 18240 22204 18480 22228
rect 18240 22142 18264 22204
rect 18456 22142 18480 22204
rect 18240 21988 18480 22142
rect 22240 22204 22480 22228
rect 22240 22142 22264 22204
rect 22456 22142 22480 22204
rect 22240 21988 22480 22142
rect 26240 22204 26480 22228
rect 26240 22142 26264 22204
rect 26456 22142 26480 22204
rect 26240 21988 26480 22142
rect 30240 22204 30480 22228
rect 30240 22142 30264 22204
rect 30456 22142 30480 22204
rect 30240 21988 30480 22142
rect 34240 22204 34480 22228
rect 34240 22142 34264 22204
rect 34456 22142 34480 22204
rect 34240 21988 34480 22142
rect 38240 22204 38480 22228
rect 38240 22142 38264 22204
rect 38456 22142 38480 22204
rect 38240 21988 38480 22142
rect 1934 21768 2254 21822
rect 360 21524 600 21548
rect 360 21332 384 21524
rect 576 21332 600 21524
rect 1934 21528 1960 21768
rect 2182 21528 2200 21768
rect 2206 21528 2254 21768
rect 3602 21771 3690 21776
rect 3602 21693 3607 21771
rect 3685 21693 3690 21771
rect 3602 21688 3690 21693
rect 5934 21768 6254 21822
rect 1934 21502 2254 21528
rect 4360 21524 4600 21548
rect 360 21308 600 21332
rect 4360 21332 4384 21524
rect 4576 21332 4600 21524
rect 5934 21528 5960 21768
rect 6182 21528 6200 21768
rect 6206 21528 6254 21768
rect 7602 21771 7690 21776
rect 7602 21693 7607 21771
rect 7685 21693 7690 21771
rect 7602 21688 7690 21693
rect 9934 21768 10254 21822
rect 5934 21502 6254 21528
rect 8360 21524 8600 21548
rect 2810 21319 2946 21324
rect 2810 21245 2815 21319
rect 2941 21245 2946 21319
rect 4360 21308 4600 21332
rect 8360 21332 8384 21524
rect 8576 21332 8600 21524
rect 9934 21528 9960 21768
rect 10182 21528 10200 21768
rect 10206 21528 10254 21768
rect 11602 21771 11690 21776
rect 11602 21693 11607 21771
rect 11685 21693 11690 21771
rect 11602 21688 11690 21693
rect 13934 21768 14254 21822
rect 9934 21502 10254 21528
rect 12360 21524 12600 21548
rect 6810 21319 6946 21324
rect 2810 21240 2946 21245
rect 6810 21245 6815 21319
rect 6941 21245 6946 21319
rect 8360 21308 8600 21332
rect 12360 21332 12384 21524
rect 12576 21332 12600 21524
rect 13934 21528 13960 21768
rect 14182 21528 14200 21768
rect 14206 21528 14254 21768
rect 15602 21771 15690 21776
rect 15602 21693 15607 21771
rect 15685 21693 15690 21771
rect 15602 21688 15690 21693
rect 17934 21768 18254 21822
rect 13934 21502 14254 21528
rect 16360 21524 16600 21548
rect 10810 21319 10946 21324
rect 6810 21240 6946 21245
rect 10810 21245 10815 21319
rect 10941 21245 10946 21319
rect 12360 21308 12600 21332
rect 16360 21332 16384 21524
rect 16576 21332 16600 21524
rect 17934 21528 17960 21768
rect 18182 21528 18200 21768
rect 18206 21528 18254 21768
rect 19602 21771 19690 21776
rect 19602 21693 19607 21771
rect 19685 21693 19690 21771
rect 19602 21688 19690 21693
rect 21934 21768 22254 21822
rect 17934 21502 18254 21528
rect 20360 21524 20600 21548
rect 14810 21319 14946 21324
rect 10810 21240 10946 21245
rect 14810 21245 14815 21319
rect 14941 21245 14946 21319
rect 16360 21308 16600 21332
rect 20360 21332 20384 21524
rect 20576 21332 20600 21524
rect 21934 21528 21960 21768
rect 22182 21528 22200 21768
rect 22206 21528 22254 21768
rect 23602 21771 23690 21776
rect 23602 21693 23607 21771
rect 23685 21693 23690 21771
rect 23602 21688 23690 21693
rect 25934 21768 26254 21822
rect 21934 21502 22254 21528
rect 24360 21524 24600 21548
rect 18810 21319 18946 21324
rect 14810 21240 14946 21245
rect 18810 21245 18815 21319
rect 18941 21245 18946 21319
rect 20360 21308 20600 21332
rect 24360 21332 24384 21524
rect 24576 21332 24600 21524
rect 25934 21528 25960 21768
rect 26182 21528 26200 21768
rect 26206 21528 26254 21768
rect 27602 21771 27690 21776
rect 27602 21693 27607 21771
rect 27685 21693 27690 21771
rect 27602 21688 27690 21693
rect 29934 21768 30254 21822
rect 25934 21502 26254 21528
rect 28360 21524 28600 21548
rect 22810 21319 22946 21324
rect 18810 21240 18946 21245
rect 22810 21245 22815 21319
rect 22941 21245 22946 21319
rect 24360 21308 24600 21332
rect 28360 21332 28384 21524
rect 28576 21332 28600 21524
rect 29934 21528 29960 21768
rect 30182 21528 30200 21768
rect 30206 21528 30254 21768
rect 31602 21771 31690 21776
rect 31602 21693 31607 21771
rect 31685 21693 31690 21771
rect 31602 21688 31690 21693
rect 33934 21768 34254 21822
rect 29934 21502 30254 21528
rect 32360 21524 32600 21548
rect 26810 21319 26946 21324
rect 22810 21240 22946 21245
rect 26810 21245 26815 21319
rect 26941 21245 26946 21319
rect 28360 21308 28600 21332
rect 32360 21332 32384 21524
rect 32576 21332 32600 21524
rect 33934 21528 33960 21768
rect 34182 21528 34200 21768
rect 34206 21528 34254 21768
rect 35602 21771 35690 21776
rect 35602 21693 35607 21771
rect 35685 21693 35690 21771
rect 35602 21688 35690 21693
rect 37934 21768 38254 21822
rect 33934 21502 34254 21528
rect 36360 21524 36600 21548
rect 30810 21319 30946 21324
rect 26810 21240 26946 21245
rect 30810 21245 30815 21319
rect 30941 21245 30946 21319
rect 32360 21308 32600 21332
rect 36360 21332 36384 21524
rect 36576 21332 36600 21524
rect 37934 21528 37960 21768
rect 38182 21528 38200 21768
rect 38206 21528 38254 21768
rect 39602 21771 39690 21776
rect 39602 21693 39607 21771
rect 39685 21693 39690 21771
rect 39602 21688 39690 21693
rect 37934 21502 38254 21528
rect 34810 21319 34946 21324
rect 30810 21240 30946 21245
rect 34810 21245 34815 21319
rect 34941 21245 34946 21319
rect 36360 21308 36600 21332
rect 38810 21319 38946 21324
rect 34810 21240 34946 21245
rect 38810 21245 38815 21319
rect 38941 21245 38946 21319
rect 38810 21240 38946 21245
rect 2338 21181 2518 21182
rect 2338 21003 2339 21181
rect 2517 21003 2518 21181
rect 2338 21002 2518 21003
rect 6338 21181 6518 21182
rect 6338 21003 6339 21181
rect 6517 21003 6518 21181
rect 6338 21002 6518 21003
rect 10338 21181 10518 21182
rect 10338 21003 10339 21181
rect 10517 21003 10518 21181
rect 10338 21002 10518 21003
rect 14338 21181 14518 21182
rect 14338 21003 14339 21181
rect 14517 21003 14518 21181
rect 14338 21002 14518 21003
rect 18338 21181 18518 21182
rect 18338 21003 18339 21181
rect 18517 21003 18518 21181
rect 18338 21002 18518 21003
rect 22338 21181 22518 21182
rect 22338 21003 22339 21181
rect 22517 21003 22518 21181
rect 22338 21002 22518 21003
rect 26338 21181 26518 21182
rect 26338 21003 26339 21181
rect 26517 21003 26518 21181
rect 26338 21002 26518 21003
rect 30338 21181 30518 21182
rect 30338 21003 30339 21181
rect 30517 21003 30518 21181
rect 30338 21002 30518 21003
rect 34338 21181 34518 21182
rect 34338 21003 34339 21181
rect 34517 21003 34518 21181
rect 34338 21002 34518 21003
rect 38338 21181 38518 21182
rect 38338 21003 38339 21181
rect 38517 21003 38518 21181
rect 38338 21002 38518 21003
rect 390 20607 570 20608
rect 390 20429 391 20607
rect 569 20429 570 20607
rect 3734 20604 3740 20610
rect 3780 20604 3786 20610
rect 4390 20607 4570 20608
rect 3728 20598 3734 20604
rect 3786 20598 3792 20604
rect 3728 20552 3734 20558
rect 3786 20552 3792 20558
rect 3734 20546 3740 20552
rect 3780 20546 3786 20552
rect 390 20428 570 20429
rect 4390 20429 4391 20607
rect 4569 20429 4570 20607
rect 7734 20604 7740 20610
rect 7780 20604 7786 20610
rect 8390 20607 8570 20608
rect 7728 20598 7734 20604
rect 7786 20598 7792 20604
rect 7728 20552 7734 20558
rect 7786 20552 7792 20558
rect 7734 20546 7740 20552
rect 7780 20546 7786 20552
rect 4390 20428 4570 20429
rect 8390 20429 8391 20607
rect 8569 20429 8570 20607
rect 11734 20604 11740 20610
rect 11780 20604 11786 20610
rect 12390 20607 12570 20608
rect 11728 20598 11734 20604
rect 11786 20598 11792 20604
rect 11728 20552 11734 20558
rect 11786 20552 11792 20558
rect 11734 20546 11740 20552
rect 11780 20546 11786 20552
rect 8390 20428 8570 20429
rect 12390 20429 12391 20607
rect 12569 20429 12570 20607
rect 15734 20604 15740 20610
rect 15780 20604 15786 20610
rect 16390 20607 16570 20608
rect 15728 20598 15734 20604
rect 15786 20598 15792 20604
rect 15728 20552 15734 20558
rect 15786 20552 15792 20558
rect 15734 20546 15740 20552
rect 15780 20546 15786 20552
rect 12390 20428 12570 20429
rect 16390 20429 16391 20607
rect 16569 20429 16570 20607
rect 19734 20604 19740 20610
rect 19780 20604 19786 20610
rect 20390 20607 20570 20608
rect 19728 20598 19734 20604
rect 19786 20598 19792 20604
rect 19728 20552 19734 20558
rect 19786 20552 19792 20558
rect 19734 20546 19740 20552
rect 19780 20546 19786 20552
rect 16390 20428 16570 20429
rect 20390 20429 20391 20607
rect 20569 20429 20570 20607
rect 23734 20604 23740 20610
rect 23780 20604 23786 20610
rect 24390 20607 24570 20608
rect 23728 20598 23734 20604
rect 23786 20598 23792 20604
rect 23728 20552 23734 20558
rect 23786 20552 23792 20558
rect 23734 20546 23740 20552
rect 23780 20546 23786 20552
rect 20390 20428 20570 20429
rect 24390 20429 24391 20607
rect 24569 20429 24570 20607
rect 27734 20604 27740 20610
rect 27780 20604 27786 20610
rect 28390 20607 28570 20608
rect 27728 20598 27734 20604
rect 27786 20598 27792 20604
rect 27728 20552 27734 20558
rect 27786 20552 27792 20558
rect 27734 20546 27740 20552
rect 27780 20546 27786 20552
rect 24390 20428 24570 20429
rect 28390 20429 28391 20607
rect 28569 20429 28570 20607
rect 31734 20604 31740 20610
rect 31780 20604 31786 20610
rect 32390 20607 32570 20608
rect 31728 20598 31734 20604
rect 31786 20598 31792 20604
rect 31728 20552 31734 20558
rect 31786 20552 31792 20558
rect 31734 20546 31740 20552
rect 31780 20546 31786 20552
rect 28390 20428 28570 20429
rect 32390 20429 32391 20607
rect 32569 20429 32570 20607
rect 35734 20604 35740 20610
rect 35780 20604 35786 20610
rect 36390 20607 36570 20608
rect 35728 20598 35734 20604
rect 35786 20598 35792 20604
rect 35728 20552 35734 20558
rect 35786 20552 35792 20558
rect 35734 20546 35740 20552
rect 35780 20546 35786 20552
rect 32390 20428 32570 20429
rect 36390 20429 36391 20607
rect 36569 20429 36570 20607
rect 39734 20604 39740 20610
rect 39780 20604 39786 20610
rect 39728 20598 39734 20604
rect 39786 20598 39792 20604
rect 39728 20552 39734 20558
rect 39786 20552 39792 20558
rect 39734 20546 39740 20552
rect 39780 20546 39786 20552
rect 36390 20428 36570 20429
rect 3262 20416 3268 20422
rect 3308 20416 3314 20422
rect 7262 20416 7268 20422
rect 7308 20416 7314 20422
rect 11262 20416 11268 20422
rect 11308 20416 11314 20422
rect 15262 20416 15268 20422
rect 15308 20416 15314 20422
rect 19262 20416 19268 20422
rect 19308 20416 19314 20422
rect 23262 20416 23268 20422
rect 23308 20416 23314 20422
rect 27262 20416 27268 20422
rect 27308 20416 27314 20422
rect 31262 20416 31268 20422
rect 31308 20416 31314 20422
rect 35262 20416 35268 20422
rect 35308 20416 35314 20422
rect 39262 20416 39268 20422
rect 39308 20416 39314 20422
rect 3256 20410 3262 20416
rect 3314 20410 3320 20416
rect 7256 20410 7262 20416
rect 7314 20410 7320 20416
rect 11256 20410 11262 20416
rect 11314 20410 11320 20416
rect 15256 20410 15262 20416
rect 15314 20410 15320 20416
rect 19256 20410 19262 20416
rect 19314 20410 19320 20416
rect 23256 20410 23262 20416
rect 23314 20410 23320 20416
rect 27256 20410 27262 20416
rect 27314 20410 27320 20416
rect 31256 20410 31262 20416
rect 31314 20410 31320 20416
rect 35256 20410 35262 20416
rect 35314 20410 35320 20416
rect 39256 20410 39262 20416
rect 39314 20410 39320 20416
rect 3256 20364 3262 20370
rect 3314 20364 3320 20370
rect 7256 20364 7262 20370
rect 7314 20364 7320 20370
rect 11256 20364 11262 20370
rect 11314 20364 11320 20370
rect 15256 20364 15262 20370
rect 15314 20364 15320 20370
rect 19256 20364 19262 20370
rect 19314 20364 19320 20370
rect 23256 20364 23262 20370
rect 23314 20364 23320 20370
rect 27256 20364 27262 20370
rect 27314 20364 27320 20370
rect 31256 20364 31262 20370
rect 31314 20364 31320 20370
rect 35256 20364 35262 20370
rect 35314 20364 35320 20370
rect 39256 20364 39262 20370
rect 39314 20364 39320 20370
rect 3262 20358 3268 20364
rect 3308 20358 3314 20364
rect 7262 20358 7268 20364
rect 7308 20358 7314 20364
rect 11262 20358 11268 20364
rect 11308 20358 11314 20364
rect 15262 20358 15268 20364
rect 15308 20358 15314 20364
rect 19262 20358 19268 20364
rect 19308 20358 19314 20364
rect 23262 20358 23268 20364
rect 23308 20358 23314 20364
rect 27262 20358 27268 20364
rect 27308 20358 27314 20364
rect 31262 20358 31268 20364
rect 31308 20358 31314 20364
rect 35262 20358 35268 20364
rect 35308 20358 35314 20364
rect 39262 20358 39268 20364
rect 39308 20358 39314 20364
rect 2240 19904 2480 19928
rect 2240 19712 2264 19904
rect 2456 19712 2480 19904
rect 2240 19688 2480 19712
rect 6240 19904 6480 19928
rect 6240 19712 6264 19904
rect 6456 19712 6480 19904
rect 6240 19688 6480 19712
rect 10240 19904 10480 19928
rect 10240 19712 10264 19904
rect 10456 19712 10480 19904
rect 10240 19688 10480 19712
rect 14240 19904 14480 19928
rect 14240 19712 14264 19904
rect 14456 19712 14480 19904
rect 14240 19688 14480 19712
rect 18240 19904 18480 19928
rect 18240 19712 18264 19904
rect 18456 19712 18480 19904
rect 18240 19688 18480 19712
rect 22240 19904 22480 19928
rect 22240 19712 22264 19904
rect 22456 19712 22480 19904
rect 22240 19688 22480 19712
rect 26240 19904 26480 19928
rect 26240 19712 26264 19904
rect 26456 19712 26480 19904
rect 26240 19688 26480 19712
rect 30240 19904 30480 19928
rect 30240 19712 30264 19904
rect 30456 19712 30480 19904
rect 30240 19688 30480 19712
rect 34240 19904 34480 19928
rect 34240 19712 34264 19904
rect 34456 19712 34480 19904
rect 34240 19688 34480 19712
rect 38240 19904 38480 19928
rect 38240 19712 38264 19904
rect 38456 19712 38480 19904
rect 38240 19688 38480 19712
rect 2240 19204 2480 19228
rect 2240 19142 2264 19204
rect 2456 19142 2480 19204
rect 2240 18988 2480 19142
rect 6240 19204 6480 19228
rect 6240 19142 6264 19204
rect 6456 19142 6480 19204
rect 6240 18988 6480 19142
rect 10240 19204 10480 19228
rect 10240 19142 10264 19204
rect 10456 19142 10480 19204
rect 10240 18988 10480 19142
rect 14240 19204 14480 19228
rect 14240 19142 14264 19204
rect 14456 19142 14480 19204
rect 14240 18988 14480 19142
rect 18240 19204 18480 19228
rect 18240 19142 18264 19204
rect 18456 19142 18480 19204
rect 18240 18988 18480 19142
rect 22240 19204 22480 19228
rect 22240 19142 22264 19204
rect 22456 19142 22480 19204
rect 22240 18988 22480 19142
rect 26240 19204 26480 19228
rect 26240 19142 26264 19204
rect 26456 19142 26480 19204
rect 26240 18988 26480 19142
rect 30240 19204 30480 19228
rect 30240 19142 30264 19204
rect 30456 19142 30480 19204
rect 30240 18988 30480 19142
rect 34240 19204 34480 19228
rect 34240 19142 34264 19204
rect 34456 19142 34480 19204
rect 34240 18988 34480 19142
rect 38240 19204 38480 19228
rect 38240 19142 38264 19204
rect 38456 19142 38480 19204
rect 38240 18988 38480 19142
rect 1934 18768 2254 18822
rect 360 18524 600 18548
rect 360 18332 384 18524
rect 576 18332 600 18524
rect 1934 18528 1960 18768
rect 2182 18528 2200 18768
rect 2206 18528 2254 18768
rect 3602 18771 3690 18776
rect 3602 18693 3607 18771
rect 3685 18693 3690 18771
rect 3602 18688 3690 18693
rect 5934 18768 6254 18822
rect 1934 18502 2254 18528
rect 4360 18524 4600 18548
rect 360 18308 600 18332
rect 4360 18332 4384 18524
rect 4576 18332 4600 18524
rect 5934 18528 5960 18768
rect 6182 18528 6200 18768
rect 6206 18528 6254 18768
rect 7602 18771 7690 18776
rect 7602 18693 7607 18771
rect 7685 18693 7690 18771
rect 7602 18688 7690 18693
rect 9934 18768 10254 18822
rect 5934 18502 6254 18528
rect 8360 18524 8600 18548
rect 2810 18319 2946 18324
rect 2810 18245 2815 18319
rect 2941 18245 2946 18319
rect 4360 18308 4600 18332
rect 8360 18332 8384 18524
rect 8576 18332 8600 18524
rect 9934 18528 9960 18768
rect 10182 18528 10200 18768
rect 10206 18528 10254 18768
rect 11602 18771 11690 18776
rect 11602 18693 11607 18771
rect 11685 18693 11690 18771
rect 11602 18688 11690 18693
rect 13934 18768 14254 18822
rect 9934 18502 10254 18528
rect 12360 18524 12600 18548
rect 6810 18319 6946 18324
rect 2810 18240 2946 18245
rect 6810 18245 6815 18319
rect 6941 18245 6946 18319
rect 8360 18308 8600 18332
rect 12360 18332 12384 18524
rect 12576 18332 12600 18524
rect 13934 18528 13960 18768
rect 14182 18528 14200 18768
rect 14206 18528 14254 18768
rect 15602 18771 15690 18776
rect 15602 18693 15607 18771
rect 15685 18693 15690 18771
rect 15602 18688 15690 18693
rect 17934 18768 18254 18822
rect 13934 18502 14254 18528
rect 16360 18524 16600 18548
rect 10810 18319 10946 18324
rect 6810 18240 6946 18245
rect 10810 18245 10815 18319
rect 10941 18245 10946 18319
rect 12360 18308 12600 18332
rect 16360 18332 16384 18524
rect 16576 18332 16600 18524
rect 17934 18528 17960 18768
rect 18182 18528 18200 18768
rect 18206 18528 18254 18768
rect 19602 18771 19690 18776
rect 19602 18693 19607 18771
rect 19685 18693 19690 18771
rect 19602 18688 19690 18693
rect 21934 18768 22254 18822
rect 17934 18502 18254 18528
rect 20360 18524 20600 18548
rect 14810 18319 14946 18324
rect 10810 18240 10946 18245
rect 14810 18245 14815 18319
rect 14941 18245 14946 18319
rect 16360 18308 16600 18332
rect 20360 18332 20384 18524
rect 20576 18332 20600 18524
rect 21934 18528 21960 18768
rect 22182 18528 22200 18768
rect 22206 18528 22254 18768
rect 23602 18771 23690 18776
rect 23602 18693 23607 18771
rect 23685 18693 23690 18771
rect 23602 18688 23690 18693
rect 25934 18768 26254 18822
rect 21934 18502 22254 18528
rect 24360 18524 24600 18548
rect 18810 18319 18946 18324
rect 14810 18240 14946 18245
rect 18810 18245 18815 18319
rect 18941 18245 18946 18319
rect 20360 18308 20600 18332
rect 24360 18332 24384 18524
rect 24576 18332 24600 18524
rect 25934 18528 25960 18768
rect 26182 18528 26200 18768
rect 26206 18528 26254 18768
rect 27602 18771 27690 18776
rect 27602 18693 27607 18771
rect 27685 18693 27690 18771
rect 27602 18688 27690 18693
rect 29934 18768 30254 18822
rect 25934 18502 26254 18528
rect 28360 18524 28600 18548
rect 22810 18319 22946 18324
rect 18810 18240 18946 18245
rect 22810 18245 22815 18319
rect 22941 18245 22946 18319
rect 24360 18308 24600 18332
rect 28360 18332 28384 18524
rect 28576 18332 28600 18524
rect 29934 18528 29960 18768
rect 30182 18528 30200 18768
rect 30206 18528 30254 18768
rect 31602 18771 31690 18776
rect 31602 18693 31607 18771
rect 31685 18693 31690 18771
rect 31602 18688 31690 18693
rect 33934 18768 34254 18822
rect 29934 18502 30254 18528
rect 32360 18524 32600 18548
rect 26810 18319 26946 18324
rect 22810 18240 22946 18245
rect 26810 18245 26815 18319
rect 26941 18245 26946 18319
rect 28360 18308 28600 18332
rect 32360 18332 32384 18524
rect 32576 18332 32600 18524
rect 33934 18528 33960 18768
rect 34182 18528 34200 18768
rect 34206 18528 34254 18768
rect 35602 18771 35690 18776
rect 35602 18693 35607 18771
rect 35685 18693 35690 18771
rect 35602 18688 35690 18693
rect 37934 18768 38254 18822
rect 33934 18502 34254 18528
rect 36360 18524 36600 18548
rect 30810 18319 30946 18324
rect 26810 18240 26946 18245
rect 30810 18245 30815 18319
rect 30941 18245 30946 18319
rect 32360 18308 32600 18332
rect 36360 18332 36384 18524
rect 36576 18332 36600 18524
rect 37934 18528 37960 18768
rect 38182 18528 38200 18768
rect 38206 18528 38254 18768
rect 39602 18771 39690 18776
rect 39602 18693 39607 18771
rect 39685 18693 39690 18771
rect 39602 18688 39690 18693
rect 37934 18502 38254 18528
rect 34810 18319 34946 18324
rect 30810 18240 30946 18245
rect 34810 18245 34815 18319
rect 34941 18245 34946 18319
rect 36360 18308 36600 18332
rect 38810 18319 38946 18324
rect 34810 18240 34946 18245
rect 38810 18245 38815 18319
rect 38941 18245 38946 18319
rect 38810 18240 38946 18245
rect 2338 18181 2518 18182
rect 2338 18003 2339 18181
rect 2517 18003 2518 18181
rect 2338 18002 2518 18003
rect 6338 18181 6518 18182
rect 6338 18003 6339 18181
rect 6517 18003 6518 18181
rect 6338 18002 6518 18003
rect 10338 18181 10518 18182
rect 10338 18003 10339 18181
rect 10517 18003 10518 18181
rect 10338 18002 10518 18003
rect 14338 18181 14518 18182
rect 14338 18003 14339 18181
rect 14517 18003 14518 18181
rect 14338 18002 14518 18003
rect 18338 18181 18518 18182
rect 18338 18003 18339 18181
rect 18517 18003 18518 18181
rect 18338 18002 18518 18003
rect 22338 18181 22518 18182
rect 22338 18003 22339 18181
rect 22517 18003 22518 18181
rect 22338 18002 22518 18003
rect 26338 18181 26518 18182
rect 26338 18003 26339 18181
rect 26517 18003 26518 18181
rect 26338 18002 26518 18003
rect 30338 18181 30518 18182
rect 30338 18003 30339 18181
rect 30517 18003 30518 18181
rect 30338 18002 30518 18003
rect 34338 18181 34518 18182
rect 34338 18003 34339 18181
rect 34517 18003 34518 18181
rect 34338 18002 34518 18003
rect 38338 18181 38518 18182
rect 38338 18003 38339 18181
rect 38517 18003 38518 18181
rect 38338 18002 38518 18003
rect 390 17607 570 17608
rect 390 17429 391 17607
rect 569 17429 570 17607
rect 3734 17604 3740 17610
rect 3780 17604 3786 17610
rect 4390 17607 4570 17608
rect 3728 17598 3734 17604
rect 3786 17598 3792 17604
rect 3728 17552 3734 17558
rect 3786 17552 3792 17558
rect 3734 17546 3740 17552
rect 3780 17546 3786 17552
rect 390 17428 570 17429
rect 4390 17429 4391 17607
rect 4569 17429 4570 17607
rect 7734 17604 7740 17610
rect 7780 17604 7786 17610
rect 8390 17607 8570 17608
rect 7728 17598 7734 17604
rect 7786 17598 7792 17604
rect 7728 17552 7734 17558
rect 7786 17552 7792 17558
rect 7734 17546 7740 17552
rect 7780 17546 7786 17552
rect 4390 17428 4570 17429
rect 8390 17429 8391 17607
rect 8569 17429 8570 17607
rect 11734 17604 11740 17610
rect 11780 17604 11786 17610
rect 12390 17607 12570 17608
rect 11728 17598 11734 17604
rect 11786 17598 11792 17604
rect 11728 17552 11734 17558
rect 11786 17552 11792 17558
rect 11734 17546 11740 17552
rect 11780 17546 11786 17552
rect 8390 17428 8570 17429
rect 12390 17429 12391 17607
rect 12569 17429 12570 17607
rect 15734 17604 15740 17610
rect 15780 17604 15786 17610
rect 16390 17607 16570 17608
rect 15728 17598 15734 17604
rect 15786 17598 15792 17604
rect 15728 17552 15734 17558
rect 15786 17552 15792 17558
rect 15734 17546 15740 17552
rect 15780 17546 15786 17552
rect 12390 17428 12570 17429
rect 16390 17429 16391 17607
rect 16569 17429 16570 17607
rect 19734 17604 19740 17610
rect 19780 17604 19786 17610
rect 20390 17607 20570 17608
rect 19728 17598 19734 17604
rect 19786 17598 19792 17604
rect 19728 17552 19734 17558
rect 19786 17552 19792 17558
rect 19734 17546 19740 17552
rect 19780 17546 19786 17552
rect 16390 17428 16570 17429
rect 20390 17429 20391 17607
rect 20569 17429 20570 17607
rect 23734 17604 23740 17610
rect 23780 17604 23786 17610
rect 24390 17607 24570 17608
rect 23728 17598 23734 17604
rect 23786 17598 23792 17604
rect 23728 17552 23734 17558
rect 23786 17552 23792 17558
rect 23734 17546 23740 17552
rect 23780 17546 23786 17552
rect 20390 17428 20570 17429
rect 24390 17429 24391 17607
rect 24569 17429 24570 17607
rect 27734 17604 27740 17610
rect 27780 17604 27786 17610
rect 28390 17607 28570 17608
rect 27728 17598 27734 17604
rect 27786 17598 27792 17604
rect 27728 17552 27734 17558
rect 27786 17552 27792 17558
rect 27734 17546 27740 17552
rect 27780 17546 27786 17552
rect 24390 17428 24570 17429
rect 28390 17429 28391 17607
rect 28569 17429 28570 17607
rect 31734 17604 31740 17610
rect 31780 17604 31786 17610
rect 32390 17607 32570 17608
rect 31728 17598 31734 17604
rect 31786 17598 31792 17604
rect 31728 17552 31734 17558
rect 31786 17552 31792 17558
rect 31734 17546 31740 17552
rect 31780 17546 31786 17552
rect 28390 17428 28570 17429
rect 32390 17429 32391 17607
rect 32569 17429 32570 17607
rect 35734 17604 35740 17610
rect 35780 17604 35786 17610
rect 36390 17607 36570 17608
rect 35728 17598 35734 17604
rect 35786 17598 35792 17604
rect 35728 17552 35734 17558
rect 35786 17552 35792 17558
rect 35734 17546 35740 17552
rect 35780 17546 35786 17552
rect 32390 17428 32570 17429
rect 36390 17429 36391 17607
rect 36569 17429 36570 17607
rect 39734 17604 39740 17610
rect 39780 17604 39786 17610
rect 39728 17598 39734 17604
rect 39786 17598 39792 17604
rect 39728 17552 39734 17558
rect 39786 17552 39792 17558
rect 39734 17546 39740 17552
rect 39780 17546 39786 17552
rect 36390 17428 36570 17429
rect 3262 17416 3268 17422
rect 3308 17416 3314 17422
rect 7262 17416 7268 17422
rect 7308 17416 7314 17422
rect 11262 17416 11268 17422
rect 11308 17416 11314 17422
rect 15262 17416 15268 17422
rect 15308 17416 15314 17422
rect 19262 17416 19268 17422
rect 19308 17416 19314 17422
rect 23262 17416 23268 17422
rect 23308 17416 23314 17422
rect 27262 17416 27268 17422
rect 27308 17416 27314 17422
rect 31262 17416 31268 17422
rect 31308 17416 31314 17422
rect 35262 17416 35268 17422
rect 35308 17416 35314 17422
rect 39262 17416 39268 17422
rect 39308 17416 39314 17422
rect 3256 17410 3262 17416
rect 3314 17410 3320 17416
rect 7256 17410 7262 17416
rect 7314 17410 7320 17416
rect 11256 17410 11262 17416
rect 11314 17410 11320 17416
rect 15256 17410 15262 17416
rect 15314 17410 15320 17416
rect 19256 17410 19262 17416
rect 19314 17410 19320 17416
rect 23256 17410 23262 17416
rect 23314 17410 23320 17416
rect 27256 17410 27262 17416
rect 27314 17410 27320 17416
rect 31256 17410 31262 17416
rect 31314 17410 31320 17416
rect 35256 17410 35262 17416
rect 35314 17410 35320 17416
rect 39256 17410 39262 17416
rect 39314 17410 39320 17416
rect 3256 17364 3262 17370
rect 3314 17364 3320 17370
rect 7256 17364 7262 17370
rect 7314 17364 7320 17370
rect 11256 17364 11262 17370
rect 11314 17364 11320 17370
rect 15256 17364 15262 17370
rect 15314 17364 15320 17370
rect 19256 17364 19262 17370
rect 19314 17364 19320 17370
rect 23256 17364 23262 17370
rect 23314 17364 23320 17370
rect 27256 17364 27262 17370
rect 27314 17364 27320 17370
rect 31256 17364 31262 17370
rect 31314 17364 31320 17370
rect 35256 17364 35262 17370
rect 35314 17364 35320 17370
rect 39256 17364 39262 17370
rect 39314 17364 39320 17370
rect 3262 17358 3268 17364
rect 3308 17358 3314 17364
rect 7262 17358 7268 17364
rect 7308 17358 7314 17364
rect 11262 17358 11268 17364
rect 11308 17358 11314 17364
rect 15262 17358 15268 17364
rect 15308 17358 15314 17364
rect 19262 17358 19268 17364
rect 19308 17358 19314 17364
rect 23262 17358 23268 17364
rect 23308 17358 23314 17364
rect 27262 17358 27268 17364
rect 27308 17358 27314 17364
rect 31262 17358 31268 17364
rect 31308 17358 31314 17364
rect 35262 17358 35268 17364
rect 35308 17358 35314 17364
rect 39262 17358 39268 17364
rect 39308 17358 39314 17364
rect 2240 16904 2480 16928
rect 2240 16712 2264 16904
rect 2456 16712 2480 16904
rect 2240 16688 2480 16712
rect 6240 16904 6480 16928
rect 6240 16712 6264 16904
rect 6456 16712 6480 16904
rect 6240 16688 6480 16712
rect 10240 16904 10480 16928
rect 10240 16712 10264 16904
rect 10456 16712 10480 16904
rect 10240 16688 10480 16712
rect 14240 16904 14480 16928
rect 14240 16712 14264 16904
rect 14456 16712 14480 16904
rect 14240 16688 14480 16712
rect 18240 16904 18480 16928
rect 18240 16712 18264 16904
rect 18456 16712 18480 16904
rect 18240 16688 18480 16712
rect 22240 16904 22480 16928
rect 22240 16712 22264 16904
rect 22456 16712 22480 16904
rect 22240 16688 22480 16712
rect 26240 16904 26480 16928
rect 26240 16712 26264 16904
rect 26456 16712 26480 16904
rect 26240 16688 26480 16712
rect 30240 16904 30480 16928
rect 30240 16712 30264 16904
rect 30456 16712 30480 16904
rect 30240 16688 30480 16712
rect 34240 16904 34480 16928
rect 34240 16712 34264 16904
rect 34456 16712 34480 16904
rect 34240 16688 34480 16712
rect 38240 16904 38480 16928
rect 38240 16712 38264 16904
rect 38456 16712 38480 16904
rect 38240 16688 38480 16712
rect 2240 16204 2480 16228
rect 2240 16142 2264 16204
rect 2456 16142 2480 16204
rect 2240 15988 2480 16142
rect 6240 16204 6480 16228
rect 6240 16142 6264 16204
rect 6456 16142 6480 16204
rect 6240 15988 6480 16142
rect 10240 16204 10480 16228
rect 10240 16142 10264 16204
rect 10456 16142 10480 16204
rect 10240 15988 10480 16142
rect 14240 16204 14480 16228
rect 14240 16142 14264 16204
rect 14456 16142 14480 16204
rect 14240 15988 14480 16142
rect 18240 16204 18480 16228
rect 18240 16142 18264 16204
rect 18456 16142 18480 16204
rect 18240 15988 18480 16142
rect 22240 16204 22480 16228
rect 22240 16142 22264 16204
rect 22456 16142 22480 16204
rect 22240 15988 22480 16142
rect 26240 16204 26480 16228
rect 26240 16142 26264 16204
rect 26456 16142 26480 16204
rect 26240 15988 26480 16142
rect 30240 16204 30480 16228
rect 30240 16142 30264 16204
rect 30456 16142 30480 16204
rect 30240 15988 30480 16142
rect 34240 16204 34480 16228
rect 34240 16142 34264 16204
rect 34456 16142 34480 16204
rect 34240 15988 34480 16142
rect 38240 16204 38480 16228
rect 38240 16142 38264 16204
rect 38456 16142 38480 16204
rect 38240 15988 38480 16142
rect 1934 15768 2254 15822
rect 360 15524 600 15548
rect 360 15332 384 15524
rect 576 15332 600 15524
rect 1934 15528 1960 15768
rect 2182 15528 2200 15768
rect 2206 15528 2254 15768
rect 3602 15771 3690 15776
rect 3602 15693 3607 15771
rect 3685 15693 3690 15771
rect 3602 15688 3690 15693
rect 5934 15768 6254 15822
rect 1934 15502 2254 15528
rect 4360 15524 4600 15548
rect 360 15308 600 15332
rect 4360 15332 4384 15524
rect 4576 15332 4600 15524
rect 5934 15528 5960 15768
rect 6182 15528 6200 15768
rect 6206 15528 6254 15768
rect 7602 15771 7690 15776
rect 7602 15693 7607 15771
rect 7685 15693 7690 15771
rect 7602 15688 7690 15693
rect 9934 15768 10254 15822
rect 5934 15502 6254 15528
rect 8360 15524 8600 15548
rect 2810 15319 2946 15324
rect 2810 15245 2815 15319
rect 2941 15245 2946 15319
rect 4360 15308 4600 15332
rect 8360 15332 8384 15524
rect 8576 15332 8600 15524
rect 9934 15528 9960 15768
rect 10182 15528 10200 15768
rect 10206 15528 10254 15768
rect 11602 15771 11690 15776
rect 11602 15693 11607 15771
rect 11685 15693 11690 15771
rect 11602 15688 11690 15693
rect 13934 15768 14254 15822
rect 9934 15502 10254 15528
rect 12360 15524 12600 15548
rect 6810 15319 6946 15324
rect 2810 15240 2946 15245
rect 6810 15245 6815 15319
rect 6941 15245 6946 15319
rect 8360 15308 8600 15332
rect 12360 15332 12384 15524
rect 12576 15332 12600 15524
rect 13934 15528 13960 15768
rect 14182 15528 14200 15768
rect 14206 15528 14254 15768
rect 15602 15771 15690 15776
rect 15602 15693 15607 15771
rect 15685 15693 15690 15771
rect 15602 15688 15690 15693
rect 17934 15768 18254 15822
rect 13934 15502 14254 15528
rect 16360 15524 16600 15548
rect 10810 15319 10946 15324
rect 6810 15240 6946 15245
rect 10810 15245 10815 15319
rect 10941 15245 10946 15319
rect 12360 15308 12600 15332
rect 16360 15332 16384 15524
rect 16576 15332 16600 15524
rect 17934 15528 17960 15768
rect 18182 15528 18200 15768
rect 18206 15528 18254 15768
rect 19602 15771 19690 15776
rect 19602 15693 19607 15771
rect 19685 15693 19690 15771
rect 19602 15688 19690 15693
rect 21934 15768 22254 15822
rect 17934 15502 18254 15528
rect 20360 15524 20600 15548
rect 14810 15319 14946 15324
rect 10810 15240 10946 15245
rect 14810 15245 14815 15319
rect 14941 15245 14946 15319
rect 16360 15308 16600 15332
rect 20360 15332 20384 15524
rect 20576 15332 20600 15524
rect 21934 15528 21960 15768
rect 22182 15528 22200 15768
rect 22206 15528 22254 15768
rect 23602 15771 23690 15776
rect 23602 15693 23607 15771
rect 23685 15693 23690 15771
rect 23602 15688 23690 15693
rect 25934 15768 26254 15822
rect 21934 15502 22254 15528
rect 24360 15524 24600 15548
rect 18810 15319 18946 15324
rect 14810 15240 14946 15245
rect 18810 15245 18815 15319
rect 18941 15245 18946 15319
rect 20360 15308 20600 15332
rect 24360 15332 24384 15524
rect 24576 15332 24600 15524
rect 25934 15528 25960 15768
rect 26182 15528 26200 15768
rect 26206 15528 26254 15768
rect 27602 15771 27690 15776
rect 27602 15693 27607 15771
rect 27685 15693 27690 15771
rect 27602 15688 27690 15693
rect 29934 15768 30254 15822
rect 25934 15502 26254 15528
rect 28360 15524 28600 15548
rect 22810 15319 22946 15324
rect 18810 15240 18946 15245
rect 22810 15245 22815 15319
rect 22941 15245 22946 15319
rect 24360 15308 24600 15332
rect 28360 15332 28384 15524
rect 28576 15332 28600 15524
rect 29934 15528 29960 15768
rect 30182 15528 30200 15768
rect 30206 15528 30254 15768
rect 31602 15771 31690 15776
rect 31602 15693 31607 15771
rect 31685 15693 31690 15771
rect 31602 15688 31690 15693
rect 33934 15768 34254 15822
rect 29934 15502 30254 15528
rect 32360 15524 32600 15548
rect 26810 15319 26946 15324
rect 22810 15240 22946 15245
rect 26810 15245 26815 15319
rect 26941 15245 26946 15319
rect 28360 15308 28600 15332
rect 32360 15332 32384 15524
rect 32576 15332 32600 15524
rect 33934 15528 33960 15768
rect 34182 15528 34200 15768
rect 34206 15528 34254 15768
rect 35602 15771 35690 15776
rect 35602 15693 35607 15771
rect 35685 15693 35690 15771
rect 35602 15688 35690 15693
rect 37934 15768 38254 15822
rect 33934 15502 34254 15528
rect 36360 15524 36600 15548
rect 30810 15319 30946 15324
rect 26810 15240 26946 15245
rect 30810 15245 30815 15319
rect 30941 15245 30946 15319
rect 32360 15308 32600 15332
rect 36360 15332 36384 15524
rect 36576 15332 36600 15524
rect 37934 15528 37960 15768
rect 38182 15528 38200 15768
rect 38206 15528 38254 15768
rect 39602 15771 39690 15776
rect 39602 15693 39607 15771
rect 39685 15693 39690 15771
rect 39602 15688 39690 15693
rect 37934 15502 38254 15528
rect 34810 15319 34946 15324
rect 30810 15240 30946 15245
rect 34810 15245 34815 15319
rect 34941 15245 34946 15319
rect 36360 15308 36600 15332
rect 38810 15319 38946 15324
rect 34810 15240 34946 15245
rect 38810 15245 38815 15319
rect 38941 15245 38946 15319
rect 38810 15240 38946 15245
rect 2338 15181 2518 15182
rect 2338 15003 2339 15181
rect 2517 15003 2518 15181
rect 2338 15002 2518 15003
rect 6338 15181 6518 15182
rect 6338 15003 6339 15181
rect 6517 15003 6518 15181
rect 6338 15002 6518 15003
rect 10338 15181 10518 15182
rect 10338 15003 10339 15181
rect 10517 15003 10518 15181
rect 10338 15002 10518 15003
rect 14338 15181 14518 15182
rect 14338 15003 14339 15181
rect 14517 15003 14518 15181
rect 14338 15002 14518 15003
rect 18338 15181 18518 15182
rect 18338 15003 18339 15181
rect 18517 15003 18518 15181
rect 18338 15002 18518 15003
rect 22338 15181 22518 15182
rect 22338 15003 22339 15181
rect 22517 15003 22518 15181
rect 22338 15002 22518 15003
rect 26338 15181 26518 15182
rect 26338 15003 26339 15181
rect 26517 15003 26518 15181
rect 26338 15002 26518 15003
rect 30338 15181 30518 15182
rect 30338 15003 30339 15181
rect 30517 15003 30518 15181
rect 30338 15002 30518 15003
rect 34338 15181 34518 15182
rect 34338 15003 34339 15181
rect 34517 15003 34518 15181
rect 34338 15002 34518 15003
rect 38338 15181 38518 15182
rect 38338 15003 38339 15181
rect 38517 15003 38518 15181
rect 38338 15002 38518 15003
rect 390 14607 570 14608
rect 390 14429 391 14607
rect 569 14429 570 14607
rect 3734 14604 3740 14610
rect 3780 14604 3786 14610
rect 4390 14607 4570 14608
rect 3728 14598 3734 14604
rect 3786 14598 3792 14604
rect 3728 14552 3734 14558
rect 3786 14552 3792 14558
rect 3734 14546 3740 14552
rect 3780 14546 3786 14552
rect 390 14428 570 14429
rect 4390 14429 4391 14607
rect 4569 14429 4570 14607
rect 7734 14604 7740 14610
rect 7780 14604 7786 14610
rect 8390 14607 8570 14608
rect 7728 14598 7734 14604
rect 7786 14598 7792 14604
rect 7728 14552 7734 14558
rect 7786 14552 7792 14558
rect 7734 14546 7740 14552
rect 7780 14546 7786 14552
rect 4390 14428 4570 14429
rect 8390 14429 8391 14607
rect 8569 14429 8570 14607
rect 11734 14604 11740 14610
rect 11780 14604 11786 14610
rect 12390 14607 12570 14608
rect 11728 14598 11734 14604
rect 11786 14598 11792 14604
rect 11728 14552 11734 14558
rect 11786 14552 11792 14558
rect 11734 14546 11740 14552
rect 11780 14546 11786 14552
rect 8390 14428 8570 14429
rect 12390 14429 12391 14607
rect 12569 14429 12570 14607
rect 15734 14604 15740 14610
rect 15780 14604 15786 14610
rect 16390 14607 16570 14608
rect 15728 14598 15734 14604
rect 15786 14598 15792 14604
rect 15728 14552 15734 14558
rect 15786 14552 15792 14558
rect 15734 14546 15740 14552
rect 15780 14546 15786 14552
rect 12390 14428 12570 14429
rect 16390 14429 16391 14607
rect 16569 14429 16570 14607
rect 19734 14604 19740 14610
rect 19780 14604 19786 14610
rect 20390 14607 20570 14608
rect 19728 14598 19734 14604
rect 19786 14598 19792 14604
rect 19728 14552 19734 14558
rect 19786 14552 19792 14558
rect 19734 14546 19740 14552
rect 19780 14546 19786 14552
rect 16390 14428 16570 14429
rect 20390 14429 20391 14607
rect 20569 14429 20570 14607
rect 23734 14604 23740 14610
rect 23780 14604 23786 14610
rect 24390 14607 24570 14608
rect 23728 14598 23734 14604
rect 23786 14598 23792 14604
rect 23728 14552 23734 14558
rect 23786 14552 23792 14558
rect 23734 14546 23740 14552
rect 23780 14546 23786 14552
rect 20390 14428 20570 14429
rect 24390 14429 24391 14607
rect 24569 14429 24570 14607
rect 27734 14604 27740 14610
rect 27780 14604 27786 14610
rect 28390 14607 28570 14608
rect 27728 14598 27734 14604
rect 27786 14598 27792 14604
rect 27728 14552 27734 14558
rect 27786 14552 27792 14558
rect 27734 14546 27740 14552
rect 27780 14546 27786 14552
rect 24390 14428 24570 14429
rect 28390 14429 28391 14607
rect 28569 14429 28570 14607
rect 31734 14604 31740 14610
rect 31780 14604 31786 14610
rect 32390 14607 32570 14608
rect 31728 14598 31734 14604
rect 31786 14598 31792 14604
rect 31728 14552 31734 14558
rect 31786 14552 31792 14558
rect 31734 14546 31740 14552
rect 31780 14546 31786 14552
rect 28390 14428 28570 14429
rect 32390 14429 32391 14607
rect 32569 14429 32570 14607
rect 35734 14604 35740 14610
rect 35780 14604 35786 14610
rect 36390 14607 36570 14608
rect 35728 14598 35734 14604
rect 35786 14598 35792 14604
rect 35728 14552 35734 14558
rect 35786 14552 35792 14558
rect 35734 14546 35740 14552
rect 35780 14546 35786 14552
rect 32390 14428 32570 14429
rect 36390 14429 36391 14607
rect 36569 14429 36570 14607
rect 39734 14604 39740 14610
rect 39780 14604 39786 14610
rect 39728 14598 39734 14604
rect 39786 14598 39792 14604
rect 39728 14552 39734 14558
rect 39786 14552 39792 14558
rect 39734 14546 39740 14552
rect 39780 14546 39786 14552
rect 36390 14428 36570 14429
rect 3262 14416 3268 14422
rect 3308 14416 3314 14422
rect 7262 14416 7268 14422
rect 7308 14416 7314 14422
rect 11262 14416 11268 14422
rect 11308 14416 11314 14422
rect 15262 14416 15268 14422
rect 15308 14416 15314 14422
rect 19262 14416 19268 14422
rect 19308 14416 19314 14422
rect 23262 14416 23268 14422
rect 23308 14416 23314 14422
rect 27262 14416 27268 14422
rect 27308 14416 27314 14422
rect 31262 14416 31268 14422
rect 31308 14416 31314 14422
rect 35262 14416 35268 14422
rect 35308 14416 35314 14422
rect 39262 14416 39268 14422
rect 39308 14416 39314 14422
rect 3256 14410 3262 14416
rect 3314 14410 3320 14416
rect 7256 14410 7262 14416
rect 7314 14410 7320 14416
rect 11256 14410 11262 14416
rect 11314 14410 11320 14416
rect 15256 14410 15262 14416
rect 15314 14410 15320 14416
rect 19256 14410 19262 14416
rect 19314 14410 19320 14416
rect 23256 14410 23262 14416
rect 23314 14410 23320 14416
rect 27256 14410 27262 14416
rect 27314 14410 27320 14416
rect 31256 14410 31262 14416
rect 31314 14410 31320 14416
rect 35256 14410 35262 14416
rect 35314 14410 35320 14416
rect 39256 14410 39262 14416
rect 39314 14410 39320 14416
rect 3256 14364 3262 14370
rect 3314 14364 3320 14370
rect 7256 14364 7262 14370
rect 7314 14364 7320 14370
rect 11256 14364 11262 14370
rect 11314 14364 11320 14370
rect 15256 14364 15262 14370
rect 15314 14364 15320 14370
rect 19256 14364 19262 14370
rect 19314 14364 19320 14370
rect 23256 14364 23262 14370
rect 23314 14364 23320 14370
rect 27256 14364 27262 14370
rect 27314 14364 27320 14370
rect 31256 14364 31262 14370
rect 31314 14364 31320 14370
rect 35256 14364 35262 14370
rect 35314 14364 35320 14370
rect 39256 14364 39262 14370
rect 39314 14364 39320 14370
rect 3262 14358 3268 14364
rect 3308 14358 3314 14364
rect 7262 14358 7268 14364
rect 7308 14358 7314 14364
rect 11262 14358 11268 14364
rect 11308 14358 11314 14364
rect 15262 14358 15268 14364
rect 15308 14358 15314 14364
rect 19262 14358 19268 14364
rect 19308 14358 19314 14364
rect 23262 14358 23268 14364
rect 23308 14358 23314 14364
rect 27262 14358 27268 14364
rect 27308 14358 27314 14364
rect 31262 14358 31268 14364
rect 31308 14358 31314 14364
rect 35262 14358 35268 14364
rect 35308 14358 35314 14364
rect 39262 14358 39268 14364
rect 39308 14358 39314 14364
rect 2240 13904 2480 13928
rect 2240 13712 2264 13904
rect 2456 13712 2480 13904
rect 2240 13688 2480 13712
rect 6240 13904 6480 13928
rect 6240 13712 6264 13904
rect 6456 13712 6480 13904
rect 6240 13688 6480 13712
rect 10240 13904 10480 13928
rect 10240 13712 10264 13904
rect 10456 13712 10480 13904
rect 10240 13688 10480 13712
rect 14240 13904 14480 13928
rect 14240 13712 14264 13904
rect 14456 13712 14480 13904
rect 14240 13688 14480 13712
rect 18240 13904 18480 13928
rect 18240 13712 18264 13904
rect 18456 13712 18480 13904
rect 18240 13688 18480 13712
rect 22240 13904 22480 13928
rect 22240 13712 22264 13904
rect 22456 13712 22480 13904
rect 22240 13688 22480 13712
rect 26240 13904 26480 13928
rect 26240 13712 26264 13904
rect 26456 13712 26480 13904
rect 26240 13688 26480 13712
rect 30240 13904 30480 13928
rect 30240 13712 30264 13904
rect 30456 13712 30480 13904
rect 30240 13688 30480 13712
rect 34240 13904 34480 13928
rect 34240 13712 34264 13904
rect 34456 13712 34480 13904
rect 34240 13688 34480 13712
rect 38240 13904 38480 13928
rect 38240 13712 38264 13904
rect 38456 13712 38480 13904
rect 38240 13688 38480 13712
rect 2240 13204 2480 13228
rect 2240 13142 2264 13204
rect 2456 13142 2480 13204
rect 2240 12988 2480 13142
rect 6240 13204 6480 13228
rect 6240 13142 6264 13204
rect 6456 13142 6480 13204
rect 6240 12988 6480 13142
rect 10240 13204 10480 13228
rect 10240 13142 10264 13204
rect 10456 13142 10480 13204
rect 10240 12988 10480 13142
rect 14240 13204 14480 13228
rect 14240 13142 14264 13204
rect 14456 13142 14480 13204
rect 14240 12988 14480 13142
rect 18240 13204 18480 13228
rect 18240 13142 18264 13204
rect 18456 13142 18480 13204
rect 18240 12988 18480 13142
rect 22240 13204 22480 13228
rect 22240 13142 22264 13204
rect 22456 13142 22480 13204
rect 22240 12988 22480 13142
rect 26240 13204 26480 13228
rect 26240 13142 26264 13204
rect 26456 13142 26480 13204
rect 26240 12988 26480 13142
rect 30240 13204 30480 13228
rect 30240 13142 30264 13204
rect 30456 13142 30480 13204
rect 30240 12988 30480 13142
rect 34240 13204 34480 13228
rect 34240 13142 34264 13204
rect 34456 13142 34480 13204
rect 34240 12988 34480 13142
rect 38240 13204 38480 13228
rect 38240 13142 38264 13204
rect 38456 13142 38480 13204
rect 38240 12988 38480 13142
rect 1934 12768 2254 12822
rect 360 12524 600 12548
rect 360 12332 384 12524
rect 576 12332 600 12524
rect 1934 12528 1960 12768
rect 2182 12528 2200 12768
rect 2206 12528 2254 12768
rect 3602 12771 3690 12776
rect 3602 12693 3607 12771
rect 3685 12693 3690 12771
rect 3602 12688 3690 12693
rect 5934 12768 6254 12822
rect 1934 12502 2254 12528
rect 4360 12524 4600 12548
rect 360 12308 600 12332
rect 4360 12332 4384 12524
rect 4576 12332 4600 12524
rect 5934 12528 5960 12768
rect 6182 12528 6200 12768
rect 6206 12528 6254 12768
rect 7602 12771 7690 12776
rect 7602 12693 7607 12771
rect 7685 12693 7690 12771
rect 7602 12688 7690 12693
rect 9934 12768 10254 12822
rect 5934 12502 6254 12528
rect 8360 12524 8600 12548
rect 2810 12319 2946 12324
rect 2810 12245 2815 12319
rect 2941 12245 2946 12319
rect 4360 12308 4600 12332
rect 8360 12332 8384 12524
rect 8576 12332 8600 12524
rect 9934 12528 9960 12768
rect 10182 12528 10200 12768
rect 10206 12528 10254 12768
rect 11602 12771 11690 12776
rect 11602 12693 11607 12771
rect 11685 12693 11690 12771
rect 11602 12688 11690 12693
rect 13934 12768 14254 12822
rect 9934 12502 10254 12528
rect 12360 12524 12600 12548
rect 6810 12319 6946 12324
rect 2810 12240 2946 12245
rect 6810 12245 6815 12319
rect 6941 12245 6946 12319
rect 8360 12308 8600 12332
rect 12360 12332 12384 12524
rect 12576 12332 12600 12524
rect 13934 12528 13960 12768
rect 14182 12528 14200 12768
rect 14206 12528 14254 12768
rect 15602 12771 15690 12776
rect 15602 12693 15607 12771
rect 15685 12693 15690 12771
rect 15602 12688 15690 12693
rect 17934 12768 18254 12822
rect 13934 12502 14254 12528
rect 16360 12524 16600 12548
rect 10810 12319 10946 12324
rect 6810 12240 6946 12245
rect 10810 12245 10815 12319
rect 10941 12245 10946 12319
rect 12360 12308 12600 12332
rect 16360 12332 16384 12524
rect 16576 12332 16600 12524
rect 17934 12528 17960 12768
rect 18182 12528 18200 12768
rect 18206 12528 18254 12768
rect 19602 12771 19690 12776
rect 19602 12693 19607 12771
rect 19685 12693 19690 12771
rect 19602 12688 19690 12693
rect 21934 12768 22254 12822
rect 17934 12502 18254 12528
rect 20360 12524 20600 12548
rect 14810 12319 14946 12324
rect 10810 12240 10946 12245
rect 14810 12245 14815 12319
rect 14941 12245 14946 12319
rect 16360 12308 16600 12332
rect 20360 12332 20384 12524
rect 20576 12332 20600 12524
rect 21934 12528 21960 12768
rect 22182 12528 22200 12768
rect 22206 12528 22254 12768
rect 23602 12771 23690 12776
rect 23602 12693 23607 12771
rect 23685 12693 23690 12771
rect 23602 12688 23690 12693
rect 25934 12768 26254 12822
rect 21934 12502 22254 12528
rect 24360 12524 24600 12548
rect 18810 12319 18946 12324
rect 14810 12240 14946 12245
rect 18810 12245 18815 12319
rect 18941 12245 18946 12319
rect 20360 12308 20600 12332
rect 24360 12332 24384 12524
rect 24576 12332 24600 12524
rect 25934 12528 25960 12768
rect 26182 12528 26200 12768
rect 26206 12528 26254 12768
rect 27602 12771 27690 12776
rect 27602 12693 27607 12771
rect 27685 12693 27690 12771
rect 27602 12688 27690 12693
rect 29934 12768 30254 12822
rect 25934 12502 26254 12528
rect 28360 12524 28600 12548
rect 22810 12319 22946 12324
rect 18810 12240 18946 12245
rect 22810 12245 22815 12319
rect 22941 12245 22946 12319
rect 24360 12308 24600 12332
rect 28360 12332 28384 12524
rect 28576 12332 28600 12524
rect 29934 12528 29960 12768
rect 30182 12528 30200 12768
rect 30206 12528 30254 12768
rect 31602 12771 31690 12776
rect 31602 12693 31607 12771
rect 31685 12693 31690 12771
rect 31602 12688 31690 12693
rect 33934 12768 34254 12822
rect 29934 12502 30254 12528
rect 32360 12524 32600 12548
rect 26810 12319 26946 12324
rect 22810 12240 22946 12245
rect 26810 12245 26815 12319
rect 26941 12245 26946 12319
rect 28360 12308 28600 12332
rect 32360 12332 32384 12524
rect 32576 12332 32600 12524
rect 33934 12528 33960 12768
rect 34182 12528 34200 12768
rect 34206 12528 34254 12768
rect 35602 12771 35690 12776
rect 35602 12693 35607 12771
rect 35685 12693 35690 12771
rect 35602 12688 35690 12693
rect 37934 12768 38254 12822
rect 33934 12502 34254 12528
rect 36360 12524 36600 12548
rect 30810 12319 30946 12324
rect 26810 12240 26946 12245
rect 30810 12245 30815 12319
rect 30941 12245 30946 12319
rect 32360 12308 32600 12332
rect 36360 12332 36384 12524
rect 36576 12332 36600 12524
rect 37934 12528 37960 12768
rect 38182 12528 38200 12768
rect 38206 12528 38254 12768
rect 39602 12771 39690 12776
rect 39602 12693 39607 12771
rect 39685 12693 39690 12771
rect 39602 12688 39690 12693
rect 37934 12502 38254 12528
rect 34810 12319 34946 12324
rect 30810 12240 30946 12245
rect 34810 12245 34815 12319
rect 34941 12245 34946 12319
rect 36360 12308 36600 12332
rect 38810 12319 38946 12324
rect 34810 12240 34946 12245
rect 38810 12245 38815 12319
rect 38941 12245 38946 12319
rect 38810 12240 38946 12245
rect 2338 12181 2518 12182
rect 2338 12003 2339 12181
rect 2517 12003 2518 12181
rect 2338 12002 2518 12003
rect 6338 12181 6518 12182
rect 6338 12003 6339 12181
rect 6517 12003 6518 12181
rect 6338 12002 6518 12003
rect 10338 12181 10518 12182
rect 10338 12003 10339 12181
rect 10517 12003 10518 12181
rect 10338 12002 10518 12003
rect 14338 12181 14518 12182
rect 14338 12003 14339 12181
rect 14517 12003 14518 12181
rect 14338 12002 14518 12003
rect 18338 12181 18518 12182
rect 18338 12003 18339 12181
rect 18517 12003 18518 12181
rect 18338 12002 18518 12003
rect 22338 12181 22518 12182
rect 22338 12003 22339 12181
rect 22517 12003 22518 12181
rect 22338 12002 22518 12003
rect 26338 12181 26518 12182
rect 26338 12003 26339 12181
rect 26517 12003 26518 12181
rect 26338 12002 26518 12003
rect 30338 12181 30518 12182
rect 30338 12003 30339 12181
rect 30517 12003 30518 12181
rect 30338 12002 30518 12003
rect 34338 12181 34518 12182
rect 34338 12003 34339 12181
rect 34517 12003 34518 12181
rect 34338 12002 34518 12003
rect 38338 12181 38518 12182
rect 38338 12003 38339 12181
rect 38517 12003 38518 12181
rect 38338 12002 38518 12003
rect 390 11607 570 11608
rect 390 11429 391 11607
rect 569 11429 570 11607
rect 3734 11604 3740 11610
rect 3780 11604 3786 11610
rect 4390 11607 4570 11608
rect 3728 11598 3734 11604
rect 3786 11598 3792 11604
rect 3728 11552 3734 11558
rect 3786 11552 3792 11558
rect 3734 11546 3740 11552
rect 3780 11546 3786 11552
rect 390 11428 570 11429
rect 4390 11429 4391 11607
rect 4569 11429 4570 11607
rect 7734 11604 7740 11610
rect 7780 11604 7786 11610
rect 8390 11607 8570 11608
rect 7728 11598 7734 11604
rect 7786 11598 7792 11604
rect 7728 11552 7734 11558
rect 7786 11552 7792 11558
rect 7734 11546 7740 11552
rect 7780 11546 7786 11552
rect 4390 11428 4570 11429
rect 8390 11429 8391 11607
rect 8569 11429 8570 11607
rect 11734 11604 11740 11610
rect 11780 11604 11786 11610
rect 12390 11607 12570 11608
rect 11728 11598 11734 11604
rect 11786 11598 11792 11604
rect 11728 11552 11734 11558
rect 11786 11552 11792 11558
rect 11734 11546 11740 11552
rect 11780 11546 11786 11552
rect 8390 11428 8570 11429
rect 12390 11429 12391 11607
rect 12569 11429 12570 11607
rect 15734 11604 15740 11610
rect 15780 11604 15786 11610
rect 16390 11607 16570 11608
rect 15728 11598 15734 11604
rect 15786 11598 15792 11604
rect 15728 11552 15734 11558
rect 15786 11552 15792 11558
rect 15734 11546 15740 11552
rect 15780 11546 15786 11552
rect 12390 11428 12570 11429
rect 16390 11429 16391 11607
rect 16569 11429 16570 11607
rect 19734 11604 19740 11610
rect 19780 11604 19786 11610
rect 20390 11607 20570 11608
rect 19728 11598 19734 11604
rect 19786 11598 19792 11604
rect 19728 11552 19734 11558
rect 19786 11552 19792 11558
rect 19734 11546 19740 11552
rect 19780 11546 19786 11552
rect 16390 11428 16570 11429
rect 20390 11429 20391 11607
rect 20569 11429 20570 11607
rect 23734 11604 23740 11610
rect 23780 11604 23786 11610
rect 24390 11607 24570 11608
rect 23728 11598 23734 11604
rect 23786 11598 23792 11604
rect 23728 11552 23734 11558
rect 23786 11552 23792 11558
rect 23734 11546 23740 11552
rect 23780 11546 23786 11552
rect 20390 11428 20570 11429
rect 24390 11429 24391 11607
rect 24569 11429 24570 11607
rect 27734 11604 27740 11610
rect 27780 11604 27786 11610
rect 28390 11607 28570 11608
rect 27728 11598 27734 11604
rect 27786 11598 27792 11604
rect 27728 11552 27734 11558
rect 27786 11552 27792 11558
rect 27734 11546 27740 11552
rect 27780 11546 27786 11552
rect 24390 11428 24570 11429
rect 28390 11429 28391 11607
rect 28569 11429 28570 11607
rect 31734 11604 31740 11610
rect 31780 11604 31786 11610
rect 32390 11607 32570 11608
rect 31728 11598 31734 11604
rect 31786 11598 31792 11604
rect 31728 11552 31734 11558
rect 31786 11552 31792 11558
rect 31734 11546 31740 11552
rect 31780 11546 31786 11552
rect 28390 11428 28570 11429
rect 32390 11429 32391 11607
rect 32569 11429 32570 11607
rect 35734 11604 35740 11610
rect 35780 11604 35786 11610
rect 36390 11607 36570 11608
rect 35728 11598 35734 11604
rect 35786 11598 35792 11604
rect 35728 11552 35734 11558
rect 35786 11552 35792 11558
rect 35734 11546 35740 11552
rect 35780 11546 35786 11552
rect 32390 11428 32570 11429
rect 36390 11429 36391 11607
rect 36569 11429 36570 11607
rect 39734 11604 39740 11610
rect 39780 11604 39786 11610
rect 39728 11598 39734 11604
rect 39786 11598 39792 11604
rect 39728 11552 39734 11558
rect 39786 11552 39792 11558
rect 39734 11546 39740 11552
rect 39780 11546 39786 11552
rect 36390 11428 36570 11429
rect 3262 11416 3268 11422
rect 3308 11416 3314 11422
rect 7262 11416 7268 11422
rect 7308 11416 7314 11422
rect 11262 11416 11268 11422
rect 11308 11416 11314 11422
rect 15262 11416 15268 11422
rect 15308 11416 15314 11422
rect 19262 11416 19268 11422
rect 19308 11416 19314 11422
rect 23262 11416 23268 11422
rect 23308 11416 23314 11422
rect 27262 11416 27268 11422
rect 27308 11416 27314 11422
rect 31262 11416 31268 11422
rect 31308 11416 31314 11422
rect 35262 11416 35268 11422
rect 35308 11416 35314 11422
rect 39262 11416 39268 11422
rect 39308 11416 39314 11422
rect 3256 11410 3262 11416
rect 3314 11410 3320 11416
rect 7256 11410 7262 11416
rect 7314 11410 7320 11416
rect 11256 11410 11262 11416
rect 11314 11410 11320 11416
rect 15256 11410 15262 11416
rect 15314 11410 15320 11416
rect 19256 11410 19262 11416
rect 19314 11410 19320 11416
rect 23256 11410 23262 11416
rect 23314 11410 23320 11416
rect 27256 11410 27262 11416
rect 27314 11410 27320 11416
rect 31256 11410 31262 11416
rect 31314 11410 31320 11416
rect 35256 11410 35262 11416
rect 35314 11410 35320 11416
rect 39256 11410 39262 11416
rect 39314 11410 39320 11416
rect 3256 11364 3262 11370
rect 3314 11364 3320 11370
rect 7256 11364 7262 11370
rect 7314 11364 7320 11370
rect 11256 11364 11262 11370
rect 11314 11364 11320 11370
rect 15256 11364 15262 11370
rect 15314 11364 15320 11370
rect 19256 11364 19262 11370
rect 19314 11364 19320 11370
rect 23256 11364 23262 11370
rect 23314 11364 23320 11370
rect 27256 11364 27262 11370
rect 27314 11364 27320 11370
rect 31256 11364 31262 11370
rect 31314 11364 31320 11370
rect 35256 11364 35262 11370
rect 35314 11364 35320 11370
rect 39256 11364 39262 11370
rect 39314 11364 39320 11370
rect 3262 11358 3268 11364
rect 3308 11358 3314 11364
rect 7262 11358 7268 11364
rect 7308 11358 7314 11364
rect 11262 11358 11268 11364
rect 11308 11358 11314 11364
rect 15262 11358 15268 11364
rect 15308 11358 15314 11364
rect 19262 11358 19268 11364
rect 19308 11358 19314 11364
rect 23262 11358 23268 11364
rect 23308 11358 23314 11364
rect 27262 11358 27268 11364
rect 27308 11358 27314 11364
rect 31262 11358 31268 11364
rect 31308 11358 31314 11364
rect 35262 11358 35268 11364
rect 35308 11358 35314 11364
rect 39262 11358 39268 11364
rect 39308 11358 39314 11364
rect 2240 10904 2480 10928
rect 2240 10712 2264 10904
rect 2456 10712 2480 10904
rect 2240 10688 2480 10712
rect 6240 10904 6480 10928
rect 6240 10712 6264 10904
rect 6456 10712 6480 10904
rect 6240 10688 6480 10712
rect 10240 10904 10480 10928
rect 10240 10712 10264 10904
rect 10456 10712 10480 10904
rect 10240 10688 10480 10712
rect 14240 10904 14480 10928
rect 14240 10712 14264 10904
rect 14456 10712 14480 10904
rect 14240 10688 14480 10712
rect 18240 10904 18480 10928
rect 18240 10712 18264 10904
rect 18456 10712 18480 10904
rect 18240 10688 18480 10712
rect 22240 10904 22480 10928
rect 22240 10712 22264 10904
rect 22456 10712 22480 10904
rect 22240 10688 22480 10712
rect 26240 10904 26480 10928
rect 26240 10712 26264 10904
rect 26456 10712 26480 10904
rect 26240 10688 26480 10712
rect 30240 10904 30480 10928
rect 30240 10712 30264 10904
rect 30456 10712 30480 10904
rect 30240 10688 30480 10712
rect 34240 10904 34480 10928
rect 34240 10712 34264 10904
rect 34456 10712 34480 10904
rect 34240 10688 34480 10712
rect 38240 10904 38480 10928
rect 38240 10712 38264 10904
rect 38456 10712 38480 10904
rect 38240 10688 38480 10712
rect 2240 10204 2480 10228
rect 2240 10142 2264 10204
rect 2456 10142 2480 10204
rect 2240 9988 2480 10142
rect 6240 10204 6480 10228
rect 6240 10142 6264 10204
rect 6456 10142 6480 10204
rect 6240 9988 6480 10142
rect 10240 10204 10480 10228
rect 10240 10142 10264 10204
rect 10456 10142 10480 10204
rect 10240 9988 10480 10142
rect 14240 10204 14480 10228
rect 14240 10142 14264 10204
rect 14456 10142 14480 10204
rect 14240 9988 14480 10142
rect 18240 10204 18480 10228
rect 18240 10142 18264 10204
rect 18456 10142 18480 10204
rect 18240 9988 18480 10142
rect 22240 10204 22480 10228
rect 22240 10142 22264 10204
rect 22456 10142 22480 10204
rect 22240 9988 22480 10142
rect 26240 10204 26480 10228
rect 26240 10142 26264 10204
rect 26456 10142 26480 10204
rect 26240 9988 26480 10142
rect 30240 10204 30480 10228
rect 30240 10142 30264 10204
rect 30456 10142 30480 10204
rect 30240 9988 30480 10142
rect 34240 10204 34480 10228
rect 34240 10142 34264 10204
rect 34456 10142 34480 10204
rect 34240 9988 34480 10142
rect 38240 10204 38480 10228
rect 38240 10142 38264 10204
rect 38456 10142 38480 10204
rect 38240 9988 38480 10142
rect 1934 9768 2254 9822
rect 360 9524 600 9548
rect 360 9332 384 9524
rect 576 9332 600 9524
rect 1934 9528 1960 9768
rect 2182 9528 2200 9768
rect 2206 9528 2254 9768
rect 3602 9771 3690 9776
rect 3602 9693 3607 9771
rect 3685 9693 3690 9771
rect 3602 9688 3690 9693
rect 5934 9768 6254 9822
rect 1934 9502 2254 9528
rect 4360 9524 4600 9548
rect 360 9308 600 9332
rect 4360 9332 4384 9524
rect 4576 9332 4600 9524
rect 5934 9528 5960 9768
rect 6182 9528 6200 9768
rect 6206 9528 6254 9768
rect 7602 9771 7690 9776
rect 7602 9693 7607 9771
rect 7685 9693 7690 9771
rect 7602 9688 7690 9693
rect 9934 9768 10254 9822
rect 5934 9502 6254 9528
rect 8360 9524 8600 9548
rect 2810 9319 2946 9324
rect 2810 9245 2815 9319
rect 2941 9245 2946 9319
rect 4360 9308 4600 9332
rect 8360 9332 8384 9524
rect 8576 9332 8600 9524
rect 9934 9528 9960 9768
rect 10182 9528 10200 9768
rect 10206 9528 10254 9768
rect 11602 9771 11690 9776
rect 11602 9693 11607 9771
rect 11685 9693 11690 9771
rect 11602 9688 11690 9693
rect 13934 9768 14254 9822
rect 9934 9502 10254 9528
rect 12360 9524 12600 9548
rect 6810 9319 6946 9324
rect 2810 9240 2946 9245
rect 6810 9245 6815 9319
rect 6941 9245 6946 9319
rect 8360 9308 8600 9332
rect 12360 9332 12384 9524
rect 12576 9332 12600 9524
rect 13934 9528 13960 9768
rect 14182 9528 14200 9768
rect 14206 9528 14254 9768
rect 15602 9771 15690 9776
rect 15602 9693 15607 9771
rect 15685 9693 15690 9771
rect 15602 9688 15690 9693
rect 17934 9768 18254 9822
rect 13934 9502 14254 9528
rect 16360 9524 16600 9548
rect 10810 9319 10946 9324
rect 6810 9240 6946 9245
rect 10810 9245 10815 9319
rect 10941 9245 10946 9319
rect 12360 9308 12600 9332
rect 16360 9332 16384 9524
rect 16576 9332 16600 9524
rect 17934 9528 17960 9768
rect 18182 9528 18200 9768
rect 18206 9528 18254 9768
rect 19602 9771 19690 9776
rect 19602 9693 19607 9771
rect 19685 9693 19690 9771
rect 19602 9688 19690 9693
rect 21934 9768 22254 9822
rect 17934 9502 18254 9528
rect 20360 9524 20600 9548
rect 14810 9319 14946 9324
rect 10810 9240 10946 9245
rect 14810 9245 14815 9319
rect 14941 9245 14946 9319
rect 16360 9308 16600 9332
rect 20360 9332 20384 9524
rect 20576 9332 20600 9524
rect 21934 9528 21960 9768
rect 22182 9528 22200 9768
rect 22206 9528 22254 9768
rect 23602 9771 23690 9776
rect 23602 9693 23607 9771
rect 23685 9693 23690 9771
rect 23602 9688 23690 9693
rect 25934 9768 26254 9822
rect 21934 9502 22254 9528
rect 24360 9524 24600 9548
rect 18810 9319 18946 9324
rect 14810 9240 14946 9245
rect 18810 9245 18815 9319
rect 18941 9245 18946 9319
rect 20360 9308 20600 9332
rect 24360 9332 24384 9524
rect 24576 9332 24600 9524
rect 25934 9528 25960 9768
rect 26182 9528 26200 9768
rect 26206 9528 26254 9768
rect 27602 9771 27690 9776
rect 27602 9693 27607 9771
rect 27685 9693 27690 9771
rect 27602 9688 27690 9693
rect 29934 9768 30254 9822
rect 25934 9502 26254 9528
rect 28360 9524 28600 9548
rect 22810 9319 22946 9324
rect 18810 9240 18946 9245
rect 22810 9245 22815 9319
rect 22941 9245 22946 9319
rect 24360 9308 24600 9332
rect 28360 9332 28384 9524
rect 28576 9332 28600 9524
rect 29934 9528 29960 9768
rect 30182 9528 30200 9768
rect 30206 9528 30254 9768
rect 31602 9771 31690 9776
rect 31602 9693 31607 9771
rect 31685 9693 31690 9771
rect 31602 9688 31690 9693
rect 33934 9768 34254 9822
rect 29934 9502 30254 9528
rect 32360 9524 32600 9548
rect 26810 9319 26946 9324
rect 22810 9240 22946 9245
rect 26810 9245 26815 9319
rect 26941 9245 26946 9319
rect 28360 9308 28600 9332
rect 32360 9332 32384 9524
rect 32576 9332 32600 9524
rect 33934 9528 33960 9768
rect 34182 9528 34200 9768
rect 34206 9528 34254 9768
rect 35602 9771 35690 9776
rect 35602 9693 35607 9771
rect 35685 9693 35690 9771
rect 35602 9688 35690 9693
rect 37934 9768 38254 9822
rect 33934 9502 34254 9528
rect 36360 9524 36600 9548
rect 30810 9319 30946 9324
rect 26810 9240 26946 9245
rect 30810 9245 30815 9319
rect 30941 9245 30946 9319
rect 32360 9308 32600 9332
rect 36360 9332 36384 9524
rect 36576 9332 36600 9524
rect 37934 9528 37960 9768
rect 38182 9528 38200 9768
rect 38206 9528 38254 9768
rect 39602 9771 39690 9776
rect 39602 9693 39607 9771
rect 39685 9693 39690 9771
rect 39602 9688 39690 9693
rect 37934 9502 38254 9528
rect 34810 9319 34946 9324
rect 30810 9240 30946 9245
rect 34810 9245 34815 9319
rect 34941 9245 34946 9319
rect 36360 9308 36600 9332
rect 38810 9319 38946 9324
rect 34810 9240 34946 9245
rect 38810 9245 38815 9319
rect 38941 9245 38946 9319
rect 38810 9240 38946 9245
rect 2338 9181 2518 9182
rect 2338 9003 2339 9181
rect 2517 9003 2518 9181
rect 2338 9002 2518 9003
rect 6338 9181 6518 9182
rect 6338 9003 6339 9181
rect 6517 9003 6518 9181
rect 6338 9002 6518 9003
rect 10338 9181 10518 9182
rect 10338 9003 10339 9181
rect 10517 9003 10518 9181
rect 10338 9002 10518 9003
rect 14338 9181 14518 9182
rect 14338 9003 14339 9181
rect 14517 9003 14518 9181
rect 14338 9002 14518 9003
rect 18338 9181 18518 9182
rect 18338 9003 18339 9181
rect 18517 9003 18518 9181
rect 18338 9002 18518 9003
rect 22338 9181 22518 9182
rect 22338 9003 22339 9181
rect 22517 9003 22518 9181
rect 22338 9002 22518 9003
rect 26338 9181 26518 9182
rect 26338 9003 26339 9181
rect 26517 9003 26518 9181
rect 26338 9002 26518 9003
rect 30338 9181 30518 9182
rect 30338 9003 30339 9181
rect 30517 9003 30518 9181
rect 30338 9002 30518 9003
rect 34338 9181 34518 9182
rect 34338 9003 34339 9181
rect 34517 9003 34518 9181
rect 34338 9002 34518 9003
rect 38338 9181 38518 9182
rect 38338 9003 38339 9181
rect 38517 9003 38518 9181
rect 38338 9002 38518 9003
rect 390 8607 570 8608
rect 390 8429 391 8607
rect 569 8429 570 8607
rect 3734 8604 3740 8610
rect 3780 8604 3786 8610
rect 4390 8607 4570 8608
rect 3728 8598 3734 8604
rect 3786 8598 3792 8604
rect 3728 8552 3734 8558
rect 3786 8552 3792 8558
rect 3734 8546 3740 8552
rect 3780 8546 3786 8552
rect 390 8428 570 8429
rect 4390 8429 4391 8607
rect 4569 8429 4570 8607
rect 7734 8604 7740 8610
rect 7780 8604 7786 8610
rect 8390 8607 8570 8608
rect 7728 8598 7734 8604
rect 7786 8598 7792 8604
rect 7728 8552 7734 8558
rect 7786 8552 7792 8558
rect 7734 8546 7740 8552
rect 7780 8546 7786 8552
rect 4390 8428 4570 8429
rect 8390 8429 8391 8607
rect 8569 8429 8570 8607
rect 11734 8604 11740 8610
rect 11780 8604 11786 8610
rect 12390 8607 12570 8608
rect 11728 8598 11734 8604
rect 11786 8598 11792 8604
rect 11728 8552 11734 8558
rect 11786 8552 11792 8558
rect 11734 8546 11740 8552
rect 11780 8546 11786 8552
rect 8390 8428 8570 8429
rect 12390 8429 12391 8607
rect 12569 8429 12570 8607
rect 15734 8604 15740 8610
rect 15780 8604 15786 8610
rect 16390 8607 16570 8608
rect 15728 8598 15734 8604
rect 15786 8598 15792 8604
rect 15728 8552 15734 8558
rect 15786 8552 15792 8558
rect 15734 8546 15740 8552
rect 15780 8546 15786 8552
rect 12390 8428 12570 8429
rect 16390 8429 16391 8607
rect 16569 8429 16570 8607
rect 19734 8604 19740 8610
rect 19780 8604 19786 8610
rect 20390 8607 20570 8608
rect 19728 8598 19734 8604
rect 19786 8598 19792 8604
rect 19728 8552 19734 8558
rect 19786 8552 19792 8558
rect 19734 8546 19740 8552
rect 19780 8546 19786 8552
rect 16390 8428 16570 8429
rect 20390 8429 20391 8607
rect 20569 8429 20570 8607
rect 23734 8604 23740 8610
rect 23780 8604 23786 8610
rect 24390 8607 24570 8608
rect 23728 8598 23734 8604
rect 23786 8598 23792 8604
rect 23728 8552 23734 8558
rect 23786 8552 23792 8558
rect 23734 8546 23740 8552
rect 23780 8546 23786 8552
rect 20390 8428 20570 8429
rect 24390 8429 24391 8607
rect 24569 8429 24570 8607
rect 27734 8604 27740 8610
rect 27780 8604 27786 8610
rect 28390 8607 28570 8608
rect 27728 8598 27734 8604
rect 27786 8598 27792 8604
rect 27728 8552 27734 8558
rect 27786 8552 27792 8558
rect 27734 8546 27740 8552
rect 27780 8546 27786 8552
rect 24390 8428 24570 8429
rect 28390 8429 28391 8607
rect 28569 8429 28570 8607
rect 31734 8604 31740 8610
rect 31780 8604 31786 8610
rect 32390 8607 32570 8608
rect 31728 8598 31734 8604
rect 31786 8598 31792 8604
rect 31728 8552 31734 8558
rect 31786 8552 31792 8558
rect 31734 8546 31740 8552
rect 31780 8546 31786 8552
rect 28390 8428 28570 8429
rect 32390 8429 32391 8607
rect 32569 8429 32570 8607
rect 35734 8604 35740 8610
rect 35780 8604 35786 8610
rect 36390 8607 36570 8608
rect 35728 8598 35734 8604
rect 35786 8598 35792 8604
rect 35728 8552 35734 8558
rect 35786 8552 35792 8558
rect 35734 8546 35740 8552
rect 35780 8546 35786 8552
rect 32390 8428 32570 8429
rect 36390 8429 36391 8607
rect 36569 8429 36570 8607
rect 39734 8604 39740 8610
rect 39780 8604 39786 8610
rect 39728 8598 39734 8604
rect 39786 8598 39792 8604
rect 39728 8552 39734 8558
rect 39786 8552 39792 8558
rect 39734 8546 39740 8552
rect 39780 8546 39786 8552
rect 36390 8428 36570 8429
rect 3262 8416 3268 8422
rect 3308 8416 3314 8422
rect 7262 8416 7268 8422
rect 7308 8416 7314 8422
rect 11262 8416 11268 8422
rect 11308 8416 11314 8422
rect 15262 8416 15268 8422
rect 15308 8416 15314 8422
rect 19262 8416 19268 8422
rect 19308 8416 19314 8422
rect 23262 8416 23268 8422
rect 23308 8416 23314 8422
rect 27262 8416 27268 8422
rect 27308 8416 27314 8422
rect 31262 8416 31268 8422
rect 31308 8416 31314 8422
rect 35262 8416 35268 8422
rect 35308 8416 35314 8422
rect 39262 8416 39268 8422
rect 39308 8416 39314 8422
rect 3256 8410 3262 8416
rect 3314 8410 3320 8416
rect 7256 8410 7262 8416
rect 7314 8410 7320 8416
rect 11256 8410 11262 8416
rect 11314 8410 11320 8416
rect 15256 8410 15262 8416
rect 15314 8410 15320 8416
rect 19256 8410 19262 8416
rect 19314 8410 19320 8416
rect 23256 8410 23262 8416
rect 23314 8410 23320 8416
rect 27256 8410 27262 8416
rect 27314 8410 27320 8416
rect 31256 8410 31262 8416
rect 31314 8410 31320 8416
rect 35256 8410 35262 8416
rect 35314 8410 35320 8416
rect 39256 8410 39262 8416
rect 39314 8410 39320 8416
rect 3256 8364 3262 8370
rect 3314 8364 3320 8370
rect 7256 8364 7262 8370
rect 7314 8364 7320 8370
rect 11256 8364 11262 8370
rect 11314 8364 11320 8370
rect 15256 8364 15262 8370
rect 15314 8364 15320 8370
rect 19256 8364 19262 8370
rect 19314 8364 19320 8370
rect 23256 8364 23262 8370
rect 23314 8364 23320 8370
rect 27256 8364 27262 8370
rect 27314 8364 27320 8370
rect 31256 8364 31262 8370
rect 31314 8364 31320 8370
rect 35256 8364 35262 8370
rect 35314 8364 35320 8370
rect 39256 8364 39262 8370
rect 39314 8364 39320 8370
rect 3262 8358 3268 8364
rect 3308 8358 3314 8364
rect 7262 8358 7268 8364
rect 7308 8358 7314 8364
rect 11262 8358 11268 8364
rect 11308 8358 11314 8364
rect 15262 8358 15268 8364
rect 15308 8358 15314 8364
rect 19262 8358 19268 8364
rect 19308 8358 19314 8364
rect 23262 8358 23268 8364
rect 23308 8358 23314 8364
rect 27262 8358 27268 8364
rect 27308 8358 27314 8364
rect 31262 8358 31268 8364
rect 31308 8358 31314 8364
rect 35262 8358 35268 8364
rect 35308 8358 35314 8364
rect 39262 8358 39268 8364
rect 39308 8358 39314 8364
rect 2240 7904 2480 7928
rect 2240 7712 2264 7904
rect 2456 7712 2480 7904
rect 2240 7688 2480 7712
rect 6240 7904 6480 7928
rect 6240 7712 6264 7904
rect 6456 7712 6480 7904
rect 6240 7688 6480 7712
rect 10240 7904 10480 7928
rect 10240 7712 10264 7904
rect 10456 7712 10480 7904
rect 10240 7688 10480 7712
rect 14240 7904 14480 7928
rect 14240 7712 14264 7904
rect 14456 7712 14480 7904
rect 14240 7688 14480 7712
rect 18240 7904 18480 7928
rect 18240 7712 18264 7904
rect 18456 7712 18480 7904
rect 18240 7688 18480 7712
rect 22240 7904 22480 7928
rect 22240 7712 22264 7904
rect 22456 7712 22480 7904
rect 22240 7688 22480 7712
rect 26240 7904 26480 7928
rect 26240 7712 26264 7904
rect 26456 7712 26480 7904
rect 26240 7688 26480 7712
rect 30240 7904 30480 7928
rect 30240 7712 30264 7904
rect 30456 7712 30480 7904
rect 30240 7688 30480 7712
rect 34240 7904 34480 7928
rect 34240 7712 34264 7904
rect 34456 7712 34480 7904
rect 34240 7688 34480 7712
rect 38240 7904 38480 7928
rect 38240 7712 38264 7904
rect 38456 7712 38480 7904
rect 38240 7688 38480 7712
rect 2240 7204 2480 7228
rect 2240 7142 2264 7204
rect 2456 7142 2480 7204
rect 2240 6988 2480 7142
rect 6240 7204 6480 7228
rect 6240 7142 6264 7204
rect 6456 7142 6480 7204
rect 6240 6988 6480 7142
rect 10240 7204 10480 7228
rect 10240 7142 10264 7204
rect 10456 7142 10480 7204
rect 10240 6988 10480 7142
rect 14240 7204 14480 7228
rect 14240 7142 14264 7204
rect 14456 7142 14480 7204
rect 14240 6988 14480 7142
rect 18240 7204 18480 7228
rect 18240 7142 18264 7204
rect 18456 7142 18480 7204
rect 18240 6988 18480 7142
rect 22240 7204 22480 7228
rect 22240 7142 22264 7204
rect 22456 7142 22480 7204
rect 22240 6988 22480 7142
rect 26240 7204 26480 7228
rect 26240 7142 26264 7204
rect 26456 7142 26480 7204
rect 26240 6988 26480 7142
rect 30240 7204 30480 7228
rect 30240 7142 30264 7204
rect 30456 7142 30480 7204
rect 30240 6988 30480 7142
rect 34240 7204 34480 7228
rect 34240 7142 34264 7204
rect 34456 7142 34480 7204
rect 34240 6988 34480 7142
rect 38240 7204 38480 7228
rect 38240 7142 38264 7204
rect 38456 7142 38480 7204
rect 38240 6988 38480 7142
rect 1934 6768 2254 6822
rect 360 6524 600 6548
rect 360 6332 384 6524
rect 576 6332 600 6524
rect 1934 6528 1960 6768
rect 2182 6528 2200 6768
rect 2206 6528 2254 6768
rect 3602 6771 3690 6776
rect 3602 6693 3607 6771
rect 3685 6693 3690 6771
rect 3602 6688 3690 6693
rect 5934 6768 6254 6822
rect 1934 6502 2254 6528
rect 4360 6524 4600 6548
rect 360 6308 600 6332
rect 4360 6332 4384 6524
rect 4576 6332 4600 6524
rect 5934 6528 5960 6768
rect 6182 6528 6200 6768
rect 6206 6528 6254 6768
rect 7602 6771 7690 6776
rect 7602 6693 7607 6771
rect 7685 6693 7690 6771
rect 7602 6688 7690 6693
rect 9934 6768 10254 6822
rect 5934 6502 6254 6528
rect 8360 6524 8600 6548
rect 2810 6319 2946 6324
rect 2810 6245 2815 6319
rect 2941 6245 2946 6319
rect 4360 6308 4600 6332
rect 8360 6332 8384 6524
rect 8576 6332 8600 6524
rect 9934 6528 9960 6768
rect 10182 6528 10200 6768
rect 10206 6528 10254 6768
rect 11602 6771 11690 6776
rect 11602 6693 11607 6771
rect 11685 6693 11690 6771
rect 11602 6688 11690 6693
rect 13934 6768 14254 6822
rect 9934 6502 10254 6528
rect 12360 6524 12600 6548
rect 6810 6319 6946 6324
rect 2810 6240 2946 6245
rect 6810 6245 6815 6319
rect 6941 6245 6946 6319
rect 8360 6308 8600 6332
rect 12360 6332 12384 6524
rect 12576 6332 12600 6524
rect 13934 6528 13960 6768
rect 14182 6528 14200 6768
rect 14206 6528 14254 6768
rect 15602 6771 15690 6776
rect 15602 6693 15607 6771
rect 15685 6693 15690 6771
rect 15602 6688 15690 6693
rect 17934 6768 18254 6822
rect 13934 6502 14254 6528
rect 16360 6524 16600 6548
rect 10810 6319 10946 6324
rect 6810 6240 6946 6245
rect 10810 6245 10815 6319
rect 10941 6245 10946 6319
rect 12360 6308 12600 6332
rect 16360 6332 16384 6524
rect 16576 6332 16600 6524
rect 17934 6528 17960 6768
rect 18182 6528 18200 6768
rect 18206 6528 18254 6768
rect 19602 6771 19690 6776
rect 19602 6693 19607 6771
rect 19685 6693 19690 6771
rect 19602 6688 19690 6693
rect 21934 6768 22254 6822
rect 17934 6502 18254 6528
rect 20360 6524 20600 6548
rect 14810 6319 14946 6324
rect 10810 6240 10946 6245
rect 14810 6245 14815 6319
rect 14941 6245 14946 6319
rect 16360 6308 16600 6332
rect 20360 6332 20384 6524
rect 20576 6332 20600 6524
rect 21934 6528 21960 6768
rect 22182 6528 22200 6768
rect 22206 6528 22254 6768
rect 23602 6771 23690 6776
rect 23602 6693 23607 6771
rect 23685 6693 23690 6771
rect 23602 6688 23690 6693
rect 25934 6768 26254 6822
rect 21934 6502 22254 6528
rect 24360 6524 24600 6548
rect 18810 6319 18946 6324
rect 14810 6240 14946 6245
rect 18810 6245 18815 6319
rect 18941 6245 18946 6319
rect 20360 6308 20600 6332
rect 24360 6332 24384 6524
rect 24576 6332 24600 6524
rect 25934 6528 25960 6768
rect 26182 6528 26200 6768
rect 26206 6528 26254 6768
rect 27602 6771 27690 6776
rect 27602 6693 27607 6771
rect 27685 6693 27690 6771
rect 27602 6688 27690 6693
rect 29934 6768 30254 6822
rect 25934 6502 26254 6528
rect 28360 6524 28600 6548
rect 22810 6319 22946 6324
rect 18810 6240 18946 6245
rect 22810 6245 22815 6319
rect 22941 6245 22946 6319
rect 24360 6308 24600 6332
rect 28360 6332 28384 6524
rect 28576 6332 28600 6524
rect 29934 6528 29960 6768
rect 30182 6528 30200 6768
rect 30206 6528 30254 6768
rect 31602 6771 31690 6776
rect 31602 6693 31607 6771
rect 31685 6693 31690 6771
rect 31602 6688 31690 6693
rect 33934 6768 34254 6822
rect 29934 6502 30254 6528
rect 32360 6524 32600 6548
rect 26810 6319 26946 6324
rect 22810 6240 22946 6245
rect 26810 6245 26815 6319
rect 26941 6245 26946 6319
rect 28360 6308 28600 6332
rect 32360 6332 32384 6524
rect 32576 6332 32600 6524
rect 33934 6528 33960 6768
rect 34182 6528 34200 6768
rect 34206 6528 34254 6768
rect 35602 6771 35690 6776
rect 35602 6693 35607 6771
rect 35685 6693 35690 6771
rect 35602 6688 35690 6693
rect 37934 6768 38254 6822
rect 33934 6502 34254 6528
rect 36360 6524 36600 6548
rect 30810 6319 30946 6324
rect 26810 6240 26946 6245
rect 30810 6245 30815 6319
rect 30941 6245 30946 6319
rect 32360 6308 32600 6332
rect 36360 6332 36384 6524
rect 36576 6332 36600 6524
rect 37934 6528 37960 6768
rect 38182 6528 38200 6768
rect 38206 6528 38254 6768
rect 39602 6771 39690 6776
rect 39602 6693 39607 6771
rect 39685 6693 39690 6771
rect 39602 6688 39690 6693
rect 37934 6502 38254 6528
rect 34810 6319 34946 6324
rect 30810 6240 30946 6245
rect 34810 6245 34815 6319
rect 34941 6245 34946 6319
rect 36360 6308 36600 6332
rect 38810 6319 38946 6324
rect 34810 6240 34946 6245
rect 38810 6245 38815 6319
rect 38941 6245 38946 6319
rect 38810 6240 38946 6245
rect 2338 6181 2518 6182
rect 2338 6003 2339 6181
rect 2517 6003 2518 6181
rect 2338 6002 2518 6003
rect 6338 6181 6518 6182
rect 6338 6003 6339 6181
rect 6517 6003 6518 6181
rect 6338 6002 6518 6003
rect 10338 6181 10518 6182
rect 10338 6003 10339 6181
rect 10517 6003 10518 6181
rect 10338 6002 10518 6003
rect 14338 6181 14518 6182
rect 14338 6003 14339 6181
rect 14517 6003 14518 6181
rect 14338 6002 14518 6003
rect 18338 6181 18518 6182
rect 18338 6003 18339 6181
rect 18517 6003 18518 6181
rect 18338 6002 18518 6003
rect 22338 6181 22518 6182
rect 22338 6003 22339 6181
rect 22517 6003 22518 6181
rect 22338 6002 22518 6003
rect 26338 6181 26518 6182
rect 26338 6003 26339 6181
rect 26517 6003 26518 6181
rect 26338 6002 26518 6003
rect 30338 6181 30518 6182
rect 30338 6003 30339 6181
rect 30517 6003 30518 6181
rect 30338 6002 30518 6003
rect 34338 6181 34518 6182
rect 34338 6003 34339 6181
rect 34517 6003 34518 6181
rect 34338 6002 34518 6003
rect 38338 6181 38518 6182
rect 38338 6003 38339 6181
rect 38517 6003 38518 6181
rect 38338 6002 38518 6003
rect 390 5607 570 5608
rect 390 5429 391 5607
rect 569 5429 570 5607
rect 3734 5604 3740 5610
rect 3780 5604 3786 5610
rect 4390 5607 4570 5608
rect 3728 5598 3734 5604
rect 3786 5598 3792 5604
rect 3728 5552 3734 5558
rect 3786 5552 3792 5558
rect 3734 5546 3740 5552
rect 3780 5546 3786 5552
rect 390 5428 570 5429
rect 4390 5429 4391 5607
rect 4569 5429 4570 5607
rect 7734 5604 7740 5610
rect 7780 5604 7786 5610
rect 8390 5607 8570 5608
rect 7728 5598 7734 5604
rect 7786 5598 7792 5604
rect 7728 5552 7734 5558
rect 7786 5552 7792 5558
rect 7734 5546 7740 5552
rect 7780 5546 7786 5552
rect 4390 5428 4570 5429
rect 8390 5429 8391 5607
rect 8569 5429 8570 5607
rect 11734 5604 11740 5610
rect 11780 5604 11786 5610
rect 12390 5607 12570 5608
rect 11728 5598 11734 5604
rect 11786 5598 11792 5604
rect 11728 5552 11734 5558
rect 11786 5552 11792 5558
rect 11734 5546 11740 5552
rect 11780 5546 11786 5552
rect 8390 5428 8570 5429
rect 12390 5429 12391 5607
rect 12569 5429 12570 5607
rect 15734 5604 15740 5610
rect 15780 5604 15786 5610
rect 16390 5607 16570 5608
rect 15728 5598 15734 5604
rect 15786 5598 15792 5604
rect 15728 5552 15734 5558
rect 15786 5552 15792 5558
rect 15734 5546 15740 5552
rect 15780 5546 15786 5552
rect 12390 5428 12570 5429
rect 16390 5429 16391 5607
rect 16569 5429 16570 5607
rect 19734 5604 19740 5610
rect 19780 5604 19786 5610
rect 20390 5607 20570 5608
rect 19728 5598 19734 5604
rect 19786 5598 19792 5604
rect 19728 5552 19734 5558
rect 19786 5552 19792 5558
rect 19734 5546 19740 5552
rect 19780 5546 19786 5552
rect 16390 5428 16570 5429
rect 20390 5429 20391 5607
rect 20569 5429 20570 5607
rect 23734 5604 23740 5610
rect 23780 5604 23786 5610
rect 24390 5607 24570 5608
rect 23728 5598 23734 5604
rect 23786 5598 23792 5604
rect 23728 5552 23734 5558
rect 23786 5552 23792 5558
rect 23734 5546 23740 5552
rect 23780 5546 23786 5552
rect 20390 5428 20570 5429
rect 24390 5429 24391 5607
rect 24569 5429 24570 5607
rect 27734 5604 27740 5610
rect 27780 5604 27786 5610
rect 28390 5607 28570 5608
rect 27728 5598 27734 5604
rect 27786 5598 27792 5604
rect 27728 5552 27734 5558
rect 27786 5552 27792 5558
rect 27734 5546 27740 5552
rect 27780 5546 27786 5552
rect 24390 5428 24570 5429
rect 28390 5429 28391 5607
rect 28569 5429 28570 5607
rect 31734 5604 31740 5610
rect 31780 5604 31786 5610
rect 32390 5607 32570 5608
rect 31728 5598 31734 5604
rect 31786 5598 31792 5604
rect 31728 5552 31734 5558
rect 31786 5552 31792 5558
rect 31734 5546 31740 5552
rect 31780 5546 31786 5552
rect 28390 5428 28570 5429
rect 32390 5429 32391 5607
rect 32569 5429 32570 5607
rect 35734 5604 35740 5610
rect 35780 5604 35786 5610
rect 36390 5607 36570 5608
rect 35728 5598 35734 5604
rect 35786 5598 35792 5604
rect 35728 5552 35734 5558
rect 35786 5552 35792 5558
rect 35734 5546 35740 5552
rect 35780 5546 35786 5552
rect 32390 5428 32570 5429
rect 36390 5429 36391 5607
rect 36569 5429 36570 5607
rect 39734 5604 39740 5610
rect 39780 5604 39786 5610
rect 39728 5598 39734 5604
rect 39786 5598 39792 5604
rect 39728 5552 39734 5558
rect 39786 5552 39792 5558
rect 39734 5546 39740 5552
rect 39780 5546 39786 5552
rect 36390 5428 36570 5429
rect 3262 5416 3268 5422
rect 3308 5416 3314 5422
rect 7262 5416 7268 5422
rect 7308 5416 7314 5422
rect 11262 5416 11268 5422
rect 11308 5416 11314 5422
rect 15262 5416 15268 5422
rect 15308 5416 15314 5422
rect 19262 5416 19268 5422
rect 19308 5416 19314 5422
rect 23262 5416 23268 5422
rect 23308 5416 23314 5422
rect 27262 5416 27268 5422
rect 27308 5416 27314 5422
rect 31262 5416 31268 5422
rect 31308 5416 31314 5422
rect 35262 5416 35268 5422
rect 35308 5416 35314 5422
rect 39262 5416 39268 5422
rect 39308 5416 39314 5422
rect 3256 5410 3262 5416
rect 3314 5410 3320 5416
rect 7256 5410 7262 5416
rect 7314 5410 7320 5416
rect 11256 5410 11262 5416
rect 11314 5410 11320 5416
rect 15256 5410 15262 5416
rect 15314 5410 15320 5416
rect 19256 5410 19262 5416
rect 19314 5410 19320 5416
rect 23256 5410 23262 5416
rect 23314 5410 23320 5416
rect 27256 5410 27262 5416
rect 27314 5410 27320 5416
rect 31256 5410 31262 5416
rect 31314 5410 31320 5416
rect 35256 5410 35262 5416
rect 35314 5410 35320 5416
rect 39256 5410 39262 5416
rect 39314 5410 39320 5416
rect 3256 5364 3262 5370
rect 3314 5364 3320 5370
rect 7256 5364 7262 5370
rect 7314 5364 7320 5370
rect 11256 5364 11262 5370
rect 11314 5364 11320 5370
rect 15256 5364 15262 5370
rect 15314 5364 15320 5370
rect 19256 5364 19262 5370
rect 19314 5364 19320 5370
rect 23256 5364 23262 5370
rect 23314 5364 23320 5370
rect 27256 5364 27262 5370
rect 27314 5364 27320 5370
rect 31256 5364 31262 5370
rect 31314 5364 31320 5370
rect 35256 5364 35262 5370
rect 35314 5364 35320 5370
rect 39256 5364 39262 5370
rect 39314 5364 39320 5370
rect 3262 5358 3268 5364
rect 3308 5358 3314 5364
rect 7262 5358 7268 5364
rect 7308 5358 7314 5364
rect 11262 5358 11268 5364
rect 11308 5358 11314 5364
rect 15262 5358 15268 5364
rect 15308 5358 15314 5364
rect 19262 5358 19268 5364
rect 19308 5358 19314 5364
rect 23262 5358 23268 5364
rect 23308 5358 23314 5364
rect 27262 5358 27268 5364
rect 27308 5358 27314 5364
rect 31262 5358 31268 5364
rect 31308 5358 31314 5364
rect 35262 5358 35268 5364
rect 35308 5358 35314 5364
rect 39262 5358 39268 5364
rect 39308 5358 39314 5364
rect 2240 4904 2480 4928
rect 2240 4712 2264 4904
rect 2456 4712 2480 4904
rect 2240 4688 2480 4712
rect 6240 4904 6480 4928
rect 6240 4712 6264 4904
rect 6456 4712 6480 4904
rect 6240 4688 6480 4712
rect 10240 4904 10480 4928
rect 10240 4712 10264 4904
rect 10456 4712 10480 4904
rect 10240 4688 10480 4712
rect 14240 4904 14480 4928
rect 14240 4712 14264 4904
rect 14456 4712 14480 4904
rect 14240 4688 14480 4712
rect 18240 4904 18480 4928
rect 18240 4712 18264 4904
rect 18456 4712 18480 4904
rect 18240 4688 18480 4712
rect 22240 4904 22480 4928
rect 22240 4712 22264 4904
rect 22456 4712 22480 4904
rect 22240 4688 22480 4712
rect 26240 4904 26480 4928
rect 26240 4712 26264 4904
rect 26456 4712 26480 4904
rect 26240 4688 26480 4712
rect 30240 4904 30480 4928
rect 30240 4712 30264 4904
rect 30456 4712 30480 4904
rect 30240 4688 30480 4712
rect 34240 4904 34480 4928
rect 34240 4712 34264 4904
rect 34456 4712 34480 4904
rect 34240 4688 34480 4712
rect 38240 4904 38480 4928
rect 38240 4712 38264 4904
rect 38456 4712 38480 4904
rect 38240 4688 38480 4712
rect 2240 4204 2480 4228
rect 2240 4142 2264 4204
rect 2456 4142 2480 4204
rect 2240 3988 2480 4142
rect 6240 4204 6480 4228
rect 6240 4142 6264 4204
rect 6456 4142 6480 4204
rect 6240 3988 6480 4142
rect 10240 4204 10480 4228
rect 10240 4142 10264 4204
rect 10456 4142 10480 4204
rect 10240 3988 10480 4142
rect 14240 4204 14480 4228
rect 14240 4142 14264 4204
rect 14456 4142 14480 4204
rect 14240 3988 14480 4142
rect 18240 4204 18480 4228
rect 18240 4142 18264 4204
rect 18456 4142 18480 4204
rect 18240 3988 18480 4142
rect 22240 4204 22480 4228
rect 22240 4142 22264 4204
rect 22456 4142 22480 4204
rect 22240 3988 22480 4142
rect 26240 4204 26480 4228
rect 26240 4142 26264 4204
rect 26456 4142 26480 4204
rect 26240 3988 26480 4142
rect 30240 4204 30480 4228
rect 30240 4142 30264 4204
rect 30456 4142 30480 4204
rect 30240 3988 30480 4142
rect 34240 4204 34480 4228
rect 34240 4142 34264 4204
rect 34456 4142 34480 4204
rect 34240 3988 34480 4142
rect 38240 4204 38480 4228
rect 38240 4142 38264 4204
rect 38456 4142 38480 4204
rect 38240 3988 38480 4142
rect 1934 3768 2254 3822
rect 360 3524 600 3548
rect 360 3332 384 3524
rect 576 3332 600 3524
rect 1934 3528 1960 3768
rect 2182 3528 2200 3768
rect 2206 3528 2254 3768
rect 3602 3771 3690 3776
rect 3602 3693 3607 3771
rect 3685 3693 3690 3771
rect 3602 3688 3690 3693
rect 5934 3768 6254 3822
rect 1934 3502 2254 3528
rect 4360 3524 4600 3548
rect 360 3308 600 3332
rect 4360 3332 4384 3524
rect 4576 3332 4600 3524
rect 5934 3528 5960 3768
rect 6182 3528 6200 3768
rect 6206 3528 6254 3768
rect 7602 3771 7690 3776
rect 7602 3693 7607 3771
rect 7685 3693 7690 3771
rect 7602 3688 7690 3693
rect 9934 3768 10254 3822
rect 5934 3502 6254 3528
rect 8360 3524 8600 3548
rect 2810 3319 2946 3324
rect 2810 3245 2815 3319
rect 2941 3245 2946 3319
rect 4360 3308 4600 3332
rect 8360 3332 8384 3524
rect 8576 3332 8600 3524
rect 9934 3528 9960 3768
rect 10182 3528 10200 3768
rect 10206 3528 10254 3768
rect 11602 3771 11690 3776
rect 11602 3693 11607 3771
rect 11685 3693 11690 3771
rect 11602 3688 11690 3693
rect 13934 3768 14254 3822
rect 9934 3502 10254 3528
rect 12360 3524 12600 3548
rect 6810 3319 6946 3324
rect 2810 3240 2946 3245
rect 6810 3245 6815 3319
rect 6941 3245 6946 3319
rect 8360 3308 8600 3332
rect 12360 3332 12384 3524
rect 12576 3332 12600 3524
rect 13934 3528 13960 3768
rect 14182 3528 14200 3768
rect 14206 3528 14254 3768
rect 15602 3771 15690 3776
rect 15602 3693 15607 3771
rect 15685 3693 15690 3771
rect 15602 3688 15690 3693
rect 17934 3768 18254 3822
rect 13934 3502 14254 3528
rect 16360 3524 16600 3548
rect 10810 3319 10946 3324
rect 6810 3240 6946 3245
rect 10810 3245 10815 3319
rect 10941 3245 10946 3319
rect 12360 3308 12600 3332
rect 16360 3332 16384 3524
rect 16576 3332 16600 3524
rect 17934 3528 17960 3768
rect 18182 3528 18200 3768
rect 18206 3528 18254 3768
rect 19602 3771 19690 3776
rect 19602 3693 19607 3771
rect 19685 3693 19690 3771
rect 19602 3688 19690 3693
rect 21934 3768 22254 3822
rect 17934 3502 18254 3528
rect 20360 3524 20600 3548
rect 14810 3319 14946 3324
rect 10810 3240 10946 3245
rect 14810 3245 14815 3319
rect 14941 3245 14946 3319
rect 16360 3308 16600 3332
rect 20360 3332 20384 3524
rect 20576 3332 20600 3524
rect 21934 3528 21960 3768
rect 22182 3528 22200 3768
rect 22206 3528 22254 3768
rect 23602 3771 23690 3776
rect 23602 3693 23607 3771
rect 23685 3693 23690 3771
rect 23602 3688 23690 3693
rect 25934 3768 26254 3822
rect 21934 3502 22254 3528
rect 24360 3524 24600 3548
rect 18810 3319 18946 3324
rect 14810 3240 14946 3245
rect 18810 3245 18815 3319
rect 18941 3245 18946 3319
rect 20360 3308 20600 3332
rect 24360 3332 24384 3524
rect 24576 3332 24600 3524
rect 25934 3528 25960 3768
rect 26182 3528 26200 3768
rect 26206 3528 26254 3768
rect 27602 3771 27690 3776
rect 27602 3693 27607 3771
rect 27685 3693 27690 3771
rect 27602 3688 27690 3693
rect 29934 3768 30254 3822
rect 25934 3502 26254 3528
rect 28360 3524 28600 3548
rect 22810 3319 22946 3324
rect 18810 3240 18946 3245
rect 22810 3245 22815 3319
rect 22941 3245 22946 3319
rect 24360 3308 24600 3332
rect 28360 3332 28384 3524
rect 28576 3332 28600 3524
rect 29934 3528 29960 3768
rect 30182 3528 30200 3768
rect 30206 3528 30254 3768
rect 31602 3771 31690 3776
rect 31602 3693 31607 3771
rect 31685 3693 31690 3771
rect 31602 3688 31690 3693
rect 33934 3768 34254 3822
rect 29934 3502 30254 3528
rect 32360 3524 32600 3548
rect 26810 3319 26946 3324
rect 22810 3240 22946 3245
rect 26810 3245 26815 3319
rect 26941 3245 26946 3319
rect 28360 3308 28600 3332
rect 32360 3332 32384 3524
rect 32576 3332 32600 3524
rect 33934 3528 33960 3768
rect 34182 3528 34200 3768
rect 34206 3528 34254 3768
rect 35602 3771 35690 3776
rect 35602 3693 35607 3771
rect 35685 3693 35690 3771
rect 35602 3688 35690 3693
rect 37934 3768 38254 3822
rect 33934 3502 34254 3528
rect 36360 3524 36600 3548
rect 30810 3319 30946 3324
rect 26810 3240 26946 3245
rect 30810 3245 30815 3319
rect 30941 3245 30946 3319
rect 32360 3308 32600 3332
rect 36360 3332 36384 3524
rect 36576 3332 36600 3524
rect 37934 3528 37960 3768
rect 38182 3528 38200 3768
rect 38206 3528 38254 3768
rect 39602 3771 39690 3776
rect 39602 3693 39607 3771
rect 39685 3693 39690 3771
rect 39602 3688 39690 3693
rect 37934 3502 38254 3528
rect 34810 3319 34946 3324
rect 30810 3240 30946 3245
rect 34810 3245 34815 3319
rect 34941 3245 34946 3319
rect 36360 3308 36600 3332
rect 38810 3319 38946 3324
rect 34810 3240 34946 3245
rect 38810 3245 38815 3319
rect 38941 3245 38946 3319
rect 38810 3240 38946 3245
rect 2338 3181 2518 3182
rect 2338 3003 2339 3181
rect 2517 3003 2518 3181
rect 2338 3002 2518 3003
rect 6338 3181 6518 3182
rect 6338 3003 6339 3181
rect 6517 3003 6518 3181
rect 6338 3002 6518 3003
rect 10338 3181 10518 3182
rect 10338 3003 10339 3181
rect 10517 3003 10518 3181
rect 10338 3002 10518 3003
rect 14338 3181 14518 3182
rect 14338 3003 14339 3181
rect 14517 3003 14518 3181
rect 14338 3002 14518 3003
rect 18338 3181 18518 3182
rect 18338 3003 18339 3181
rect 18517 3003 18518 3181
rect 18338 3002 18518 3003
rect 22338 3181 22518 3182
rect 22338 3003 22339 3181
rect 22517 3003 22518 3181
rect 22338 3002 22518 3003
rect 26338 3181 26518 3182
rect 26338 3003 26339 3181
rect 26517 3003 26518 3181
rect 26338 3002 26518 3003
rect 30338 3181 30518 3182
rect 30338 3003 30339 3181
rect 30517 3003 30518 3181
rect 30338 3002 30518 3003
rect 34338 3181 34518 3182
rect 34338 3003 34339 3181
rect 34517 3003 34518 3181
rect 34338 3002 34518 3003
rect 38338 3181 38518 3182
rect 38338 3003 38339 3181
rect 38517 3003 38518 3181
rect 38338 3002 38518 3003
rect 390 2607 570 2608
rect 390 2429 391 2607
rect 569 2429 570 2607
rect 3734 2604 3740 2610
rect 3780 2604 3786 2610
rect 4390 2607 4570 2608
rect 3728 2598 3734 2604
rect 3786 2598 3792 2604
rect 3728 2552 3734 2558
rect 3786 2552 3792 2558
rect 3734 2546 3740 2552
rect 3780 2546 3786 2552
rect 390 2428 570 2429
rect 4390 2429 4391 2607
rect 4569 2429 4570 2607
rect 7734 2604 7740 2610
rect 7780 2604 7786 2610
rect 8390 2607 8570 2608
rect 7728 2598 7734 2604
rect 7786 2598 7792 2604
rect 7728 2552 7734 2558
rect 7786 2552 7792 2558
rect 7734 2546 7740 2552
rect 7780 2546 7786 2552
rect 4390 2428 4570 2429
rect 8390 2429 8391 2607
rect 8569 2429 8570 2607
rect 11734 2604 11740 2610
rect 11780 2604 11786 2610
rect 12390 2607 12570 2608
rect 11728 2598 11734 2604
rect 11786 2598 11792 2604
rect 11728 2552 11734 2558
rect 11786 2552 11792 2558
rect 11734 2546 11740 2552
rect 11780 2546 11786 2552
rect 8390 2428 8570 2429
rect 12390 2429 12391 2607
rect 12569 2429 12570 2607
rect 15734 2604 15740 2610
rect 15780 2604 15786 2610
rect 16390 2607 16570 2608
rect 15728 2598 15734 2604
rect 15786 2598 15792 2604
rect 15728 2552 15734 2558
rect 15786 2552 15792 2558
rect 15734 2546 15740 2552
rect 15780 2546 15786 2552
rect 12390 2428 12570 2429
rect 16390 2429 16391 2607
rect 16569 2429 16570 2607
rect 19734 2604 19740 2610
rect 19780 2604 19786 2610
rect 20390 2607 20570 2608
rect 19728 2598 19734 2604
rect 19786 2598 19792 2604
rect 19728 2552 19734 2558
rect 19786 2552 19792 2558
rect 19734 2546 19740 2552
rect 19780 2546 19786 2552
rect 16390 2428 16570 2429
rect 20390 2429 20391 2607
rect 20569 2429 20570 2607
rect 23734 2604 23740 2610
rect 23780 2604 23786 2610
rect 24390 2607 24570 2608
rect 23728 2598 23734 2604
rect 23786 2598 23792 2604
rect 23728 2552 23734 2558
rect 23786 2552 23792 2558
rect 23734 2546 23740 2552
rect 23780 2546 23786 2552
rect 20390 2428 20570 2429
rect 24390 2429 24391 2607
rect 24569 2429 24570 2607
rect 27734 2604 27740 2610
rect 27780 2604 27786 2610
rect 28390 2607 28570 2608
rect 27728 2598 27734 2604
rect 27786 2598 27792 2604
rect 27728 2552 27734 2558
rect 27786 2552 27792 2558
rect 27734 2546 27740 2552
rect 27780 2546 27786 2552
rect 24390 2428 24570 2429
rect 28390 2429 28391 2607
rect 28569 2429 28570 2607
rect 31734 2604 31740 2610
rect 31780 2604 31786 2610
rect 32390 2607 32570 2608
rect 31728 2598 31734 2604
rect 31786 2598 31792 2604
rect 31728 2552 31734 2558
rect 31786 2552 31792 2558
rect 31734 2546 31740 2552
rect 31780 2546 31786 2552
rect 28390 2428 28570 2429
rect 32390 2429 32391 2607
rect 32569 2429 32570 2607
rect 35734 2604 35740 2610
rect 35780 2604 35786 2610
rect 36390 2607 36570 2608
rect 35728 2598 35734 2604
rect 35786 2598 35792 2604
rect 35728 2552 35734 2558
rect 35786 2552 35792 2558
rect 35734 2546 35740 2552
rect 35780 2546 35786 2552
rect 32390 2428 32570 2429
rect 36390 2429 36391 2607
rect 36569 2429 36570 2607
rect 39734 2604 39740 2610
rect 39780 2604 39786 2610
rect 39728 2598 39734 2604
rect 39786 2598 39792 2604
rect 39728 2552 39734 2558
rect 39786 2552 39792 2558
rect 39734 2546 39740 2552
rect 39780 2546 39786 2552
rect 36390 2428 36570 2429
rect 3262 2416 3268 2422
rect 3308 2416 3314 2422
rect 7262 2416 7268 2422
rect 7308 2416 7314 2422
rect 11262 2416 11268 2422
rect 11308 2416 11314 2422
rect 15262 2416 15268 2422
rect 15308 2416 15314 2422
rect 19262 2416 19268 2422
rect 19308 2416 19314 2422
rect 23262 2416 23268 2422
rect 23308 2416 23314 2422
rect 27262 2416 27268 2422
rect 27308 2416 27314 2422
rect 31262 2416 31268 2422
rect 31308 2416 31314 2422
rect 35262 2416 35268 2422
rect 35308 2416 35314 2422
rect 39262 2416 39268 2422
rect 39308 2416 39314 2422
rect 3256 2410 3262 2416
rect 3314 2410 3320 2416
rect 7256 2410 7262 2416
rect 7314 2410 7320 2416
rect 11256 2410 11262 2416
rect 11314 2410 11320 2416
rect 15256 2410 15262 2416
rect 15314 2410 15320 2416
rect 19256 2410 19262 2416
rect 19314 2410 19320 2416
rect 23256 2410 23262 2416
rect 23314 2410 23320 2416
rect 27256 2410 27262 2416
rect 27314 2410 27320 2416
rect 31256 2410 31262 2416
rect 31314 2410 31320 2416
rect 35256 2410 35262 2416
rect 35314 2410 35320 2416
rect 39256 2410 39262 2416
rect 39314 2410 39320 2416
rect 3256 2364 3262 2370
rect 3314 2364 3320 2370
rect 7256 2364 7262 2370
rect 7314 2364 7320 2370
rect 11256 2364 11262 2370
rect 11314 2364 11320 2370
rect 15256 2364 15262 2370
rect 15314 2364 15320 2370
rect 19256 2364 19262 2370
rect 19314 2364 19320 2370
rect 23256 2364 23262 2370
rect 23314 2364 23320 2370
rect 27256 2364 27262 2370
rect 27314 2364 27320 2370
rect 31256 2364 31262 2370
rect 31314 2364 31320 2370
rect 35256 2364 35262 2370
rect 35314 2364 35320 2370
rect 39256 2364 39262 2370
rect 39314 2364 39320 2370
rect 3262 2358 3268 2364
rect 3308 2358 3314 2364
rect 7262 2358 7268 2364
rect 7308 2358 7314 2364
rect 11262 2358 11268 2364
rect 11308 2358 11314 2364
rect 15262 2358 15268 2364
rect 15308 2358 15314 2364
rect 19262 2358 19268 2364
rect 19308 2358 19314 2364
rect 23262 2358 23268 2364
rect 23308 2358 23314 2364
rect 27262 2358 27268 2364
rect 27308 2358 27314 2364
rect 31262 2358 31268 2364
rect 31308 2358 31314 2364
rect 35262 2358 35268 2364
rect 35308 2358 35314 2364
rect 39262 2358 39268 2364
rect 39308 2358 39314 2364
rect 2240 1904 2480 1928
rect 2240 1712 2264 1904
rect 2456 1712 2480 1904
rect 2240 1688 2480 1712
rect 6240 1904 6480 1928
rect 6240 1712 6264 1904
rect 6456 1712 6480 1904
rect 6240 1688 6480 1712
rect 10240 1904 10480 1928
rect 10240 1712 10264 1904
rect 10456 1712 10480 1904
rect 10240 1688 10480 1712
rect 14240 1904 14480 1928
rect 14240 1712 14264 1904
rect 14456 1712 14480 1904
rect 14240 1688 14480 1712
rect 18240 1904 18480 1928
rect 18240 1712 18264 1904
rect 18456 1712 18480 1904
rect 18240 1688 18480 1712
rect 22240 1904 22480 1928
rect 22240 1712 22264 1904
rect 22456 1712 22480 1904
rect 22240 1688 22480 1712
rect 26240 1904 26480 1928
rect 26240 1712 26264 1904
rect 26456 1712 26480 1904
rect 26240 1688 26480 1712
rect 30240 1904 30480 1928
rect 30240 1712 30264 1904
rect 30456 1712 30480 1904
rect 30240 1688 30480 1712
rect 34240 1904 34480 1928
rect 34240 1712 34264 1904
rect 34456 1712 34480 1904
rect 34240 1688 34480 1712
rect 38240 1904 38480 1928
rect 38240 1712 38264 1904
rect 38456 1712 38480 1904
rect 38240 1688 38480 1712
rect 2240 1204 2480 1228
rect 2240 1142 2264 1204
rect 2456 1142 2480 1204
rect 2240 988 2480 1142
rect 6240 1204 6480 1228
rect 6240 1142 6264 1204
rect 6456 1142 6480 1204
rect 6240 988 6480 1142
rect 10240 1204 10480 1228
rect 10240 1142 10264 1204
rect 10456 1142 10480 1204
rect 10240 988 10480 1142
rect 14240 1204 14480 1228
rect 14240 1142 14264 1204
rect 14456 1142 14480 1204
rect 14240 988 14480 1142
rect 18240 1204 18480 1228
rect 18240 1142 18264 1204
rect 18456 1142 18480 1204
rect 18240 988 18480 1142
rect 22240 1204 22480 1228
rect 22240 1142 22264 1204
rect 22456 1142 22480 1204
rect 22240 988 22480 1142
rect 26240 1204 26480 1228
rect 26240 1142 26264 1204
rect 26456 1142 26480 1204
rect 26240 988 26480 1142
rect 30240 1204 30480 1228
rect 30240 1142 30264 1204
rect 30456 1142 30480 1204
rect 30240 988 30480 1142
rect 34240 1204 34480 1228
rect 34240 1142 34264 1204
rect 34456 1142 34480 1204
rect 34240 988 34480 1142
rect 38240 1204 38480 1228
rect 38240 1142 38264 1204
rect 38456 1142 38480 1204
rect 38240 988 38480 1142
rect 1934 768 2254 822
rect 360 524 600 548
rect 360 332 384 524
rect 576 332 600 524
rect 1934 528 1960 768
rect 2182 528 2200 768
rect 2206 528 2254 768
rect 3602 771 3690 776
rect 3602 693 3607 771
rect 3685 693 3690 771
rect 3602 688 3690 693
rect 5934 768 6254 822
rect 1934 502 2254 528
rect 4360 524 4600 548
rect 360 308 600 332
rect 4360 332 4384 524
rect 4576 332 4600 524
rect 5934 528 5960 768
rect 6182 528 6200 768
rect 6206 528 6254 768
rect 7602 771 7690 776
rect 7602 693 7607 771
rect 7685 693 7690 771
rect 7602 688 7690 693
rect 9934 768 10254 822
rect 5934 502 6254 528
rect 8360 524 8600 548
rect 2810 319 2946 324
rect 2810 245 2815 319
rect 2941 245 2946 319
rect 4360 308 4600 332
rect 8360 332 8384 524
rect 8576 332 8600 524
rect 9934 528 9960 768
rect 10182 528 10200 768
rect 10206 528 10254 768
rect 11602 771 11690 776
rect 11602 693 11607 771
rect 11685 693 11690 771
rect 11602 688 11690 693
rect 13934 768 14254 822
rect 9934 502 10254 528
rect 12360 524 12600 548
rect 6810 319 6946 324
rect 2810 240 2946 245
rect 6810 245 6815 319
rect 6941 245 6946 319
rect 8360 308 8600 332
rect 12360 332 12384 524
rect 12576 332 12600 524
rect 13934 528 13960 768
rect 14182 528 14200 768
rect 14206 528 14254 768
rect 15602 771 15690 776
rect 15602 693 15607 771
rect 15685 693 15690 771
rect 15602 688 15690 693
rect 17934 768 18254 822
rect 13934 502 14254 528
rect 16360 524 16600 548
rect 10810 319 10946 324
rect 6810 240 6946 245
rect 10810 245 10815 319
rect 10941 245 10946 319
rect 12360 308 12600 332
rect 16360 332 16384 524
rect 16576 332 16600 524
rect 17934 528 17960 768
rect 18182 528 18200 768
rect 18206 528 18254 768
rect 19602 771 19690 776
rect 19602 693 19607 771
rect 19685 693 19690 771
rect 19602 688 19690 693
rect 21934 768 22254 822
rect 17934 502 18254 528
rect 20360 524 20600 548
rect 14810 319 14946 324
rect 10810 240 10946 245
rect 14810 245 14815 319
rect 14941 245 14946 319
rect 16360 308 16600 332
rect 20360 332 20384 524
rect 20576 332 20600 524
rect 21934 528 21960 768
rect 22182 528 22200 768
rect 22206 528 22254 768
rect 23602 771 23690 776
rect 23602 693 23607 771
rect 23685 693 23690 771
rect 23602 688 23690 693
rect 25934 768 26254 822
rect 21934 502 22254 528
rect 24360 524 24600 548
rect 18810 319 18946 324
rect 14810 240 14946 245
rect 18810 245 18815 319
rect 18941 245 18946 319
rect 20360 308 20600 332
rect 24360 332 24384 524
rect 24576 332 24600 524
rect 25934 528 25960 768
rect 26182 528 26200 768
rect 26206 528 26254 768
rect 27602 771 27690 776
rect 27602 693 27607 771
rect 27685 693 27690 771
rect 27602 688 27690 693
rect 29934 768 30254 822
rect 25934 502 26254 528
rect 28360 524 28600 548
rect 22810 319 22946 324
rect 18810 240 18946 245
rect 22810 245 22815 319
rect 22941 245 22946 319
rect 24360 308 24600 332
rect 28360 332 28384 524
rect 28576 332 28600 524
rect 29934 528 29960 768
rect 30182 528 30200 768
rect 30206 528 30254 768
rect 31602 771 31690 776
rect 31602 693 31607 771
rect 31685 693 31690 771
rect 31602 688 31690 693
rect 33934 768 34254 822
rect 29934 502 30254 528
rect 32360 524 32600 548
rect 26810 319 26946 324
rect 22810 240 22946 245
rect 26810 245 26815 319
rect 26941 245 26946 319
rect 28360 308 28600 332
rect 32360 332 32384 524
rect 32576 332 32600 524
rect 33934 528 33960 768
rect 34182 528 34200 768
rect 34206 528 34254 768
rect 35602 771 35690 776
rect 35602 693 35607 771
rect 35685 693 35690 771
rect 35602 688 35690 693
rect 37934 768 38254 822
rect 33934 502 34254 528
rect 36360 524 36600 548
rect 30810 319 30946 324
rect 26810 240 26946 245
rect 30810 245 30815 319
rect 30941 245 30946 319
rect 32360 308 32600 332
rect 36360 332 36384 524
rect 36576 332 36600 524
rect 37934 528 37960 768
rect 38182 528 38200 768
rect 38206 528 38254 768
rect 39602 771 39690 776
rect 39602 693 39607 771
rect 39685 693 39690 771
rect 39602 688 39690 693
rect 37934 502 38254 528
rect 34810 319 34946 324
rect 30810 240 30946 245
rect 34810 245 34815 319
rect 34941 245 34946 319
rect 36360 308 36600 332
rect 38810 319 38946 324
rect 34810 240 34946 245
rect 38810 245 38815 319
rect 38941 245 38946 319
rect 38810 240 38946 245
rect 2338 181 2518 182
rect 2338 3 2339 181
rect 2517 3 2518 181
rect 2338 2 2518 3
rect 6338 181 6518 182
rect 6338 3 6339 181
rect 6517 3 6518 181
rect 6338 2 6518 3
rect 10338 181 10518 182
rect 10338 3 10339 181
rect 10517 3 10518 181
rect 10338 2 10518 3
rect 14338 181 14518 182
rect 14338 3 14339 181
rect 14517 3 14518 181
rect 14338 2 14518 3
rect 18338 181 18518 182
rect 18338 3 18339 181
rect 18517 3 18518 181
rect 18338 2 18518 3
rect 22338 181 22518 182
rect 22338 3 22339 181
rect 22517 3 22518 181
rect 22338 2 22518 3
rect 26338 181 26518 182
rect 26338 3 26339 181
rect 26517 3 26518 181
rect 26338 2 26518 3
rect 30338 181 30518 182
rect 30338 3 30339 181
rect 30517 3 30518 181
rect 30338 2 30518 3
rect 34338 181 34518 182
rect 34338 3 34339 181
rect 34517 3 34518 181
rect 34338 2 34518 3
rect 38338 181 38518 182
rect 38338 3 38339 181
rect 38517 3 38518 181
rect 38338 2 38518 3
rect 390 -393 570 -392
rect 390 -571 391 -393
rect 569 -571 570 -393
rect 3734 -396 3740 -390
rect 3780 -396 3786 -390
rect 4390 -393 4570 -392
rect 3728 -402 3734 -396
rect 3786 -402 3792 -396
rect 3728 -448 3734 -442
rect 3786 -448 3792 -442
rect 3734 -454 3740 -448
rect 3780 -454 3786 -448
rect 390 -572 570 -571
rect 4390 -571 4391 -393
rect 4569 -571 4570 -393
rect 7734 -396 7740 -390
rect 7780 -396 7786 -390
rect 8390 -393 8570 -392
rect 7728 -402 7734 -396
rect 7786 -402 7792 -396
rect 7728 -448 7734 -442
rect 7786 -448 7792 -442
rect 7734 -454 7740 -448
rect 7780 -454 7786 -448
rect 4390 -572 4570 -571
rect 8390 -571 8391 -393
rect 8569 -571 8570 -393
rect 11734 -396 11740 -390
rect 11780 -396 11786 -390
rect 12390 -393 12570 -392
rect 11728 -402 11734 -396
rect 11786 -402 11792 -396
rect 11728 -448 11734 -442
rect 11786 -448 11792 -442
rect 11734 -454 11740 -448
rect 11780 -454 11786 -448
rect 8390 -572 8570 -571
rect 12390 -571 12391 -393
rect 12569 -571 12570 -393
rect 15734 -396 15740 -390
rect 15780 -396 15786 -390
rect 16390 -393 16570 -392
rect 15728 -402 15734 -396
rect 15786 -402 15792 -396
rect 15728 -448 15734 -442
rect 15786 -448 15792 -442
rect 15734 -454 15740 -448
rect 15780 -454 15786 -448
rect 12390 -572 12570 -571
rect 16390 -571 16391 -393
rect 16569 -571 16570 -393
rect 19734 -396 19740 -390
rect 19780 -396 19786 -390
rect 20390 -393 20570 -392
rect 19728 -402 19734 -396
rect 19786 -402 19792 -396
rect 19728 -448 19734 -442
rect 19786 -448 19792 -442
rect 19734 -454 19740 -448
rect 19780 -454 19786 -448
rect 16390 -572 16570 -571
rect 20390 -571 20391 -393
rect 20569 -571 20570 -393
rect 23734 -396 23740 -390
rect 23780 -396 23786 -390
rect 24390 -393 24570 -392
rect 23728 -402 23734 -396
rect 23786 -402 23792 -396
rect 23728 -448 23734 -442
rect 23786 -448 23792 -442
rect 23734 -454 23740 -448
rect 23780 -454 23786 -448
rect 20390 -572 20570 -571
rect 24390 -571 24391 -393
rect 24569 -571 24570 -393
rect 27734 -396 27740 -390
rect 27780 -396 27786 -390
rect 28390 -393 28570 -392
rect 27728 -402 27734 -396
rect 27786 -402 27792 -396
rect 27728 -448 27734 -442
rect 27786 -448 27792 -442
rect 27734 -454 27740 -448
rect 27780 -454 27786 -448
rect 24390 -572 24570 -571
rect 28390 -571 28391 -393
rect 28569 -571 28570 -393
rect 31734 -396 31740 -390
rect 31780 -396 31786 -390
rect 32390 -393 32570 -392
rect 31728 -402 31734 -396
rect 31786 -402 31792 -396
rect 31728 -448 31734 -442
rect 31786 -448 31792 -442
rect 31734 -454 31740 -448
rect 31780 -454 31786 -448
rect 28390 -572 28570 -571
rect 32390 -571 32391 -393
rect 32569 -571 32570 -393
rect 35734 -396 35740 -390
rect 35780 -396 35786 -390
rect 36390 -393 36570 -392
rect 35728 -402 35734 -396
rect 35786 -402 35792 -396
rect 35728 -448 35734 -442
rect 35786 -448 35792 -442
rect 35734 -454 35740 -448
rect 35780 -454 35786 -448
rect 32390 -572 32570 -571
rect 36390 -571 36391 -393
rect 36569 -571 36570 -393
rect 39734 -396 39740 -390
rect 39780 -396 39786 -390
rect 39728 -402 39734 -396
rect 39786 -402 39792 -396
rect 39728 -448 39734 -442
rect 39786 -448 39792 -442
rect 39734 -454 39740 -448
rect 39780 -454 39786 -448
rect 36390 -572 36570 -571
rect 3262 -584 3268 -578
rect 3308 -584 3314 -578
rect 7262 -584 7268 -578
rect 7308 -584 7314 -578
rect 11262 -584 11268 -578
rect 11308 -584 11314 -578
rect 15262 -584 15268 -578
rect 15308 -584 15314 -578
rect 19262 -584 19268 -578
rect 19308 -584 19314 -578
rect 23262 -584 23268 -578
rect 23308 -584 23314 -578
rect 27262 -584 27268 -578
rect 27308 -584 27314 -578
rect 31262 -584 31268 -578
rect 31308 -584 31314 -578
rect 35262 -584 35268 -578
rect 35308 -584 35314 -578
rect 39262 -584 39268 -578
rect 39308 -584 39314 -578
rect 3256 -590 3262 -584
rect 3314 -590 3320 -584
rect 7256 -590 7262 -584
rect 7314 -590 7320 -584
rect 11256 -590 11262 -584
rect 11314 -590 11320 -584
rect 15256 -590 15262 -584
rect 15314 -590 15320 -584
rect 19256 -590 19262 -584
rect 19314 -590 19320 -584
rect 23256 -590 23262 -584
rect 23314 -590 23320 -584
rect 27256 -590 27262 -584
rect 27314 -590 27320 -584
rect 31256 -590 31262 -584
rect 31314 -590 31320 -584
rect 35256 -590 35262 -584
rect 35314 -590 35320 -584
rect 39256 -590 39262 -584
rect 39314 -590 39320 -584
rect 3256 -636 3262 -630
rect 3314 -636 3320 -630
rect 7256 -636 7262 -630
rect 7314 -636 7320 -630
rect 11256 -636 11262 -630
rect 11314 -636 11320 -630
rect 15256 -636 15262 -630
rect 15314 -636 15320 -630
rect 19256 -636 19262 -630
rect 19314 -636 19320 -630
rect 23256 -636 23262 -630
rect 23314 -636 23320 -630
rect 27256 -636 27262 -630
rect 27314 -636 27320 -630
rect 31256 -636 31262 -630
rect 31314 -636 31320 -630
rect 35256 -636 35262 -630
rect 35314 -636 35320 -630
rect 39256 -636 39262 -630
rect 39314 -636 39320 -630
rect 3262 -642 3268 -636
rect 3308 -642 3314 -636
rect 7262 -642 7268 -636
rect 7308 -642 7314 -636
rect 11262 -642 11268 -636
rect 11308 -642 11314 -636
rect 15262 -642 15268 -636
rect 15308 -642 15314 -636
rect 19262 -642 19268 -636
rect 19308 -642 19314 -636
rect 23262 -642 23268 -636
rect 23308 -642 23314 -636
rect 27262 -642 27268 -636
rect 27308 -642 27314 -636
rect 31262 -642 31268 -636
rect 31308 -642 31314 -636
rect 35262 -642 35268 -636
rect 35308 -642 35314 -636
rect 39262 -642 39268 -636
rect 39308 -642 39314 -636
rect 2240 -1096 2480 -1072
rect 2240 -1288 2264 -1096
rect 2456 -1288 2480 -1096
rect 2240 -1312 2480 -1288
rect 6240 -1096 6480 -1072
rect 6240 -1288 6264 -1096
rect 6456 -1288 6480 -1096
rect 6240 -1312 6480 -1288
rect 10240 -1096 10480 -1072
rect 10240 -1288 10264 -1096
rect 10456 -1288 10480 -1096
rect 10240 -1312 10480 -1288
rect 14240 -1096 14480 -1072
rect 14240 -1288 14264 -1096
rect 14456 -1288 14480 -1096
rect 14240 -1312 14480 -1288
rect 18240 -1096 18480 -1072
rect 18240 -1288 18264 -1096
rect 18456 -1288 18480 -1096
rect 18240 -1312 18480 -1288
rect 22240 -1096 22480 -1072
rect 22240 -1288 22264 -1096
rect 22456 -1288 22480 -1096
rect 22240 -1312 22480 -1288
rect 26240 -1096 26480 -1072
rect 26240 -1288 26264 -1096
rect 26456 -1288 26480 -1096
rect 26240 -1312 26480 -1288
rect 30240 -1096 30480 -1072
rect 30240 -1288 30264 -1096
rect 30456 -1288 30480 -1096
rect 30240 -1312 30480 -1288
rect 34240 -1096 34480 -1072
rect 34240 -1288 34264 -1096
rect 34456 -1288 34480 -1096
rect 34240 -1312 34480 -1288
rect 38240 -1096 38480 -1072
rect 38240 -1288 38264 -1096
rect 38456 -1288 38480 -1096
rect 38240 -1312 38480 -1288
use fgcell_amp_MiM_cap_1_1  fgcell_amp_MiM_cap_1_1_0
array 0 9 4000 0 9 3000
timestamp 1717628967
transform 1 0 -524 0 1 2806
box 524 -4198 4490 -1570
<< end >>
