magic
tech sky130A
timestamp 1717032084
<< end >>
