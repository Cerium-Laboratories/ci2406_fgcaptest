magic
tech sky130A
magscale 1 2
timestamp 1717562480
<< pwell >>
rect -4843 -3202 4843 3202
<< psubdiff >>
rect -4807 3132 -4711 3166
rect 4711 3132 4807 3166
rect -4807 3070 -4773 3132
rect 4773 3070 4807 3132
rect -4807 -3132 -4773 -3070
rect 4773 -3132 4807 -3070
rect -4807 -3166 -4711 -3132
rect 4711 -3166 4807 -3132
<< psubdiffcont >>
rect -4711 3132 4711 3166
rect -4807 -3070 -4773 3070
rect 4773 -3070 4807 3070
rect -4711 -3166 4711 -3132
<< xpolycontact >>
rect 4395 2604 4677 3036
rect -4677 -3036 -4395 -2604
<< xpolyres >>
rect -4677 2218 -4017 2500
rect -4677 -2604 -4395 2218
rect -4299 -2218 -4017 2218
rect -3921 2218 -3261 2500
rect -3921 -2218 -3639 2218
rect -4299 -2500 -3639 -2218
rect -3543 -2218 -3261 2218
rect -3165 2218 -2505 2500
rect -3165 -2218 -2883 2218
rect -3543 -2500 -2883 -2218
rect -2787 -2218 -2505 2218
rect -2409 2218 -1749 2500
rect -2409 -2218 -2127 2218
rect -2787 -2500 -2127 -2218
rect -2031 -2218 -1749 2218
rect -1653 2218 -993 2500
rect -1653 -2218 -1371 2218
rect -2031 -2500 -1371 -2218
rect -1275 -2218 -993 2218
rect -897 2218 -237 2500
rect -897 -2218 -615 2218
rect -1275 -2500 -615 -2218
rect -519 -2218 -237 2218
rect -141 2218 519 2500
rect -141 -2218 141 2218
rect -519 -2500 141 -2218
rect 237 -2218 519 2218
rect 615 2218 1275 2500
rect 615 -2218 897 2218
rect 237 -2500 897 -2218
rect 993 -2218 1275 2218
rect 1371 2218 2031 2500
rect 1371 -2218 1653 2218
rect 993 -2500 1653 -2218
rect 1749 -2218 2031 2218
rect 2127 2218 2787 2500
rect 2127 -2218 2409 2218
rect 1749 -2500 2409 -2218
rect 2505 -2218 2787 2218
rect 2883 2218 3543 2500
rect 2883 -2218 3165 2218
rect 2505 -2500 3165 -2218
rect 3261 -2218 3543 2218
rect 3639 2218 4299 2500
rect 3639 -2218 3921 2218
rect 3261 -2500 3921 -2218
rect 4017 -2218 4299 2218
rect 4395 -2218 4677 2604
rect 4017 -2500 4677 -2218
<< locali >>
rect -4807 3132 -4711 3166
rect 4711 3132 4807 3166
rect -4807 3070 -4773 3132
rect 4773 3070 4807 3132
rect -4807 -3132 -4773 -3070
rect 4773 -3132 4807 -3070
rect -4807 -3166 -4711 -3132
rect 4711 -3166 4807 -3132
<< properties >>
string FIXED_BBOX -4790 -3149 4790 3149
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 25.0 m 1 nx 25 wmin 1.410 lmin 0.50 rho 2000 val 934.791k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
