magic
tech sky130A
timestamp 1717597221
<< nwell >>
rect 14 213 817 445
<< pwell >>
rect 14 0 817 192
<< mvnmos >>
rect 114 129 164 179
rect 193 129 243 179
rect 272 129 322 179
rect 351 129 401 179
rect 430 129 480 179
rect 509 129 559 179
rect 588 129 638 179
rect 667 129 717 179
<< mvpmos >>
rect 114 246 164 296
rect 193 246 243 296
rect 272 246 322 296
rect 351 246 401 296
rect 430 246 480 296
rect 509 246 559 296
rect 588 246 638 296
rect 667 246 717 296
<< mvndiff >>
rect 85 173 114 179
rect 85 135 91 173
rect 108 135 114 173
rect 85 129 114 135
rect 164 173 193 179
rect 164 135 170 173
rect 187 135 193 173
rect 164 129 193 135
rect 243 173 272 179
rect 243 135 249 173
rect 266 135 272 173
rect 243 129 272 135
rect 322 173 351 179
rect 322 135 328 173
rect 345 135 351 173
rect 322 129 351 135
rect 401 173 430 179
rect 401 135 407 173
rect 424 135 430 173
rect 401 129 430 135
rect 480 173 509 179
rect 480 135 486 173
rect 503 135 509 173
rect 480 129 509 135
rect 559 173 588 179
rect 559 135 565 173
rect 582 135 588 173
rect 559 129 588 135
rect 638 173 667 179
rect 638 135 644 173
rect 661 135 667 173
rect 638 129 667 135
rect 717 173 746 179
rect 717 135 723 173
rect 740 135 746 173
rect 717 129 746 135
<< mvpdiff >>
rect 85 290 114 296
rect 85 252 91 290
rect 108 252 114 290
rect 85 246 114 252
rect 164 290 193 296
rect 164 252 170 290
rect 187 252 193 290
rect 164 246 193 252
rect 243 290 272 296
rect 243 252 249 290
rect 266 252 272 290
rect 243 246 272 252
rect 322 290 351 296
rect 322 252 328 290
rect 345 252 351 290
rect 322 246 351 252
rect 401 290 430 296
rect 401 252 407 290
rect 424 252 430 290
rect 401 246 430 252
rect 480 290 509 296
rect 480 252 486 290
rect 503 252 509 290
rect 480 246 509 252
rect 559 290 588 296
rect 559 252 565 290
rect 582 252 588 290
rect 559 246 588 252
rect 638 290 667 296
rect 638 252 644 290
rect 661 252 667 290
rect 638 246 667 252
rect 717 290 746 296
rect 717 252 723 290
rect 740 252 746 290
rect 717 246 746 252
<< mvndiffc >>
rect 91 135 108 173
rect 170 135 187 173
rect 249 135 266 173
rect 328 135 345 173
rect 407 135 424 173
rect 486 135 503 173
rect 565 135 582 173
rect 644 135 661 173
rect 723 135 740 173
<< mvpdiffc >>
rect 91 252 108 290
rect 170 252 187 290
rect 249 252 266 290
rect 328 252 345 290
rect 407 252 424 290
rect 486 252 503 290
rect 565 252 582 290
rect 644 252 661 290
rect 723 252 740 290
<< mvpsubdiff >>
rect 47 41 784 47
rect 47 24 72 41
rect 759 24 784 41
rect 47 18 784 24
<< mvnsubdiff >>
rect 47 406 784 412
rect 47 389 72 406
rect 759 389 784 406
rect 47 383 784 389
<< mvpsubdiffcont >>
rect 72 24 759 41
<< mvnsubdiffcont >>
rect 72 389 759 406
<< poly >>
rect 114 337 164 345
rect 114 320 122 337
rect 156 320 164 337
rect 114 296 164 320
rect 193 337 243 345
rect 193 320 201 337
rect 235 320 243 337
rect 193 296 243 320
rect 272 337 322 345
rect 272 320 280 337
rect 314 320 322 337
rect 272 296 322 320
rect 351 337 401 345
rect 351 320 359 337
rect 393 320 401 337
rect 351 296 401 320
rect 430 337 480 345
rect 430 320 438 337
rect 472 320 480 337
rect 430 296 480 320
rect 509 337 559 345
rect 509 320 517 337
rect 551 320 559 337
rect 509 296 559 320
rect 588 337 638 345
rect 588 320 596 337
rect 630 320 638 337
rect 588 296 638 320
rect 667 337 717 345
rect 667 320 675 337
rect 709 320 717 337
rect 667 296 717 320
rect 114 233 164 246
rect 193 233 243 246
rect 272 233 322 246
rect 351 233 401 246
rect 430 233 480 246
rect 509 233 559 246
rect 588 233 638 246
rect 667 233 717 246
rect 114 179 164 192
rect 193 179 243 192
rect 272 179 322 192
rect 351 179 401 192
rect 430 179 480 192
rect 509 179 559 192
rect 588 179 638 192
rect 667 179 717 192
rect 114 110 164 129
rect 114 93 122 110
rect 156 93 164 110
rect 114 85 164 93
rect 193 110 243 129
rect 193 93 201 110
rect 235 93 243 110
rect 193 85 243 93
rect 272 110 322 129
rect 272 93 280 110
rect 314 93 322 110
rect 272 85 322 93
rect 351 110 401 129
rect 351 93 359 110
rect 393 93 401 110
rect 351 85 401 93
rect 430 110 480 129
rect 430 93 438 110
rect 472 93 480 110
rect 430 85 480 93
rect 509 110 559 129
rect 509 93 517 110
rect 551 93 559 110
rect 509 85 559 93
rect 588 110 638 129
rect 588 93 596 110
rect 630 93 638 110
rect 588 85 638 93
rect 667 110 717 129
rect 667 93 675 110
rect 709 93 717 110
rect 667 85 717 93
<< polycont >>
rect 122 320 156 337
rect 201 320 235 337
rect 280 320 314 337
rect 359 320 393 337
rect 438 320 472 337
rect 517 320 551 337
rect 596 320 630 337
rect 675 320 709 337
rect 122 93 156 110
rect 201 93 235 110
rect 280 93 314 110
rect 359 93 393 110
rect 438 93 472 110
rect 517 93 551 110
rect 596 93 630 110
rect 675 93 709 110
<< locali >>
rect 47 389 72 406
rect 759 389 784 406
rect 114 320 122 337
rect 156 320 201 337
rect 235 320 280 337
rect 314 320 359 337
rect 393 320 438 337
rect 472 320 517 337
rect 551 320 596 337
rect 630 320 675 337
rect 709 320 717 337
rect 91 290 108 298
rect 91 173 108 252
rect 91 127 108 135
rect 170 290 187 298
rect 170 173 187 252
rect 170 127 187 135
rect 249 290 266 298
rect 249 173 266 252
rect 249 127 266 135
rect 328 290 345 298
rect 328 173 345 252
rect 328 127 345 135
rect 407 290 424 298
rect 407 173 424 252
rect 407 127 424 135
rect 486 290 503 298
rect 486 173 503 252
rect 486 127 503 135
rect 565 290 582 298
rect 565 173 582 252
rect 565 127 582 135
rect 644 290 661 298
rect 644 173 661 252
rect 644 127 661 135
rect 723 290 740 298
rect 723 173 740 252
rect 723 127 740 135
rect 114 93 122 110
rect 156 93 201 110
rect 235 93 280 110
rect 314 93 359 110
rect 393 93 438 110
rect 472 93 517 110
rect 551 93 596 110
rect 630 93 675 110
rect 709 93 717 110
rect 47 24 72 41
rect 759 24 784 41
<< viali >>
rect 72 389 759 406
rect 122 320 156 337
rect 201 320 235 337
rect 280 320 314 337
rect 359 320 393 337
rect 438 320 472 337
rect 517 320 551 337
rect 596 320 630 337
rect 675 320 709 337
rect 91 252 108 290
rect 170 135 187 173
rect 249 252 266 290
rect 328 135 345 173
rect 407 252 424 290
rect 486 135 503 173
rect 565 252 582 290
rect 644 135 661 173
rect 723 252 740 290
rect 122 93 156 110
rect 201 93 235 110
rect 280 93 314 110
rect 359 93 393 110
rect 438 93 472 110
rect 517 93 551 110
rect 596 93 630 110
rect 675 93 709 110
rect 72 24 759 41
<< metal1 >>
rect 66 406 765 409
rect 66 389 72 406
rect 759 389 765 406
rect 66 386 765 389
rect 35 340 85 367
rect 35 337 717 340
rect 35 320 122 337
rect 156 320 201 337
rect 235 320 280 337
rect 314 320 359 337
rect 393 320 438 337
rect 472 320 517 337
rect 551 320 596 337
rect 630 320 675 337
rect 709 320 717 337
rect 35 317 717 320
rect 35 290 743 296
rect 35 252 91 290
rect 108 252 249 290
rect 266 252 407 290
rect 424 252 565 290
rect 582 252 723 290
rect 740 252 743 290
rect 35 246 743 252
rect 88 173 796 179
rect 88 135 170 173
rect 187 135 328 173
rect 345 135 486 173
rect 503 135 644 173
rect 661 135 796 173
rect 88 129 796 135
rect 35 110 717 113
rect 35 93 122 110
rect 156 93 201 110
rect 235 93 280 110
rect 314 93 359 110
rect 393 93 438 110
rect 472 93 517 110
rect 551 93 596 110
rect 630 93 675 110
rect 709 93 717 110
rect 35 90 717 93
rect 35 63 85 90
rect 66 41 765 44
rect 66 24 72 41
rect 759 24 765 41
rect 66 21 765 24
<< labels >>
flabel metal1 35 246 85 296 0 FreeSans 160 0 0 0 vin
port 1 nsew
flabel metal1 746 129 796 179 0 FreeSans 160 0 0 0 vout
port 2 nsew
flabel metal1 35 317 85 367 0 FreeSans 160 0 0 0 en_b
port 4 nsew
flabel metal1 35 63 85 113 0 FreeSans 160 0 0 0 en
port 3 nsew
flabel metal1 66 386 89 409 0 FreeSans 160 0 0 0 vdd
port 5 nsew
flabel metal1 66 21 89 44 0 FreeSans 160 0 0 0 vss
port 6 nsew
<< end >>
