** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/top_fgcaptest.sch
.subckt top_fgcaptest PAD_VINJ PAD_VCTRL PAD_VOUT VPWR VGND
*.PININFO PAD_VINJ:B PAD_VCTRL:I PAD_VOUT:O VPWR:I VGND:I
x1 vinj VGND net3 net4 net1 VPWR net5[9] net5[8] net5[7] net5[6] net5[5] net5[4] net5[3] net5[2] net5[1] net5[0] net6[19] net6[18]
+ net6[17] net6[16] net6[15] net6[14] net6[13] net6[12] net6[11] net6[10] net6[9] net6[8] net6[7] net6[6] net6[5] net6[4] net6[3] net6[2]
+ net6[1] net6[0] array_core
xp1 net7 vinj VGND PAD_VINJ sky130_ef_io__analog_minesd_pad_short
xp2 net1 VGND VGND PAD_VCTRL sky130_ef_io__analog_minesd_pad_short
xp3 net2 vinj VGND PAD_VOUT sky130_ef_io__analog_minesd_pad_short
.ends

* expanding   symbol:  array_core.sym # of pins=8
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core.sch
.subckt array_core vinj VGND vtun vb vctrl VPWR addr[9] addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0]
+ vout[19] vout[18] vout[17] vout[16] vout[15] vout[14] vout[13] vout[12] vout[11] vout[10] vout[9] vout[8] vout[7] vout[6] vout[5] vout[4]
+ vout[3] vout[2] vout[1] vout[0]
*.PININFO vinj:I VGND:I vtun:I vb:I vctrl:I vout[19:0]:O addr[9:0]:I VPWR:I
x1 net1 net2 net3[9] net3[8] net3[7] net3[6] net3[5] net3[4] net3[3] net3[2] net3[1] net3[0] net4[9] net4[8] net4[7] net4[6]
+ net4[5] net4[4] net4[3] net4[2] net4[1] net4[0] net5[9] net5[8] net5[7] net5[6] net5[5] net5[4] net5[3] net5[2] net5[1] net5[0] net6 net7
+ net8 net9[9] net9[8] net9[7] net9[6] net9[5] net9[4] net9[3] net9[2] net9[1] net9[0] array_core_block0
x2 net10 net11 net12[9] net12[8] net12[7] net12[6] net12[5] net12[4] net12[3] net12[2] net12[1] net12[0] net13[9] net13[8]
+ net13[7] net13[6] net13[5] net13[4] net13[3] net13[2] net13[1] net13[0] net14[9] net14[8] net14[7] net14[6] net14[5] net14[4] net14[3]
+ net14[2] net14[1] net14[0] net15 net16 net17 net18[9] net18[8] net18[7] net18[6] net18[5] net18[4] net18[3] net18[2] net18[1] net18[0]
+ array_core_block1
x3 net19 net20 net21[9] net21[8] net21[7] net21[6] net21[5] net21[4] net21[3] net21[2] net21[1] net21[0] net22[9] net22[8]
+ net22[7] net22[6] net22[5] net22[4] net22[3] net22[2] net22[1] net22[0] net23[9] net23[8] net23[7] net23[6] net23[5] net23[4] net23[3]
+ net23[2] net23[1] net23[0] net24 net25 net26 net27[9] net27[8] net27[7] net27[6] net27[5] net27[4] net27[3] net27[2] net27[1] net27[0]
+ array_core_block2
x4 net28 net29 net30[9] net30[8] net30[7] net30[6] net30[5] net30[4] net30[3] net30[2] net30[1] net30[0] net31[9] net31[8]
+ net31[7] net31[6] net31[5] net31[4] net31[3] net31[2] net31[1] net31[0] net32[9] net32[8] net32[7] net32[6] net32[5] net32[4] net32[3]
+ net32[2] net32[1] net32[0] net33 net34 net35 net36[9] net36[8] net36[7] net36[6] net36[5] net36[4] net36[3] net36[2] net36[1] net36[0]
+ array_core_block3
x5 net37 net38 net39[9] net39[8] net39[7] net39[6] net39[5] net39[4] net39[3] net39[2] net39[1] net39[0] net40[9] net40[8]
+ net40[7] net40[6] net40[5] net40[4] net40[3] net40[2] net40[1] net40[0] net41[9] net41[8] net41[7] net41[6] net41[5] net41[4] net41[3]
+ net41[2] net41[1] net41[0] net42 net43 net44 net45[9] net45[8] net45[7] net45[6] net45[5] net45[4] net45[3] net45[2] net45[1] net45[0]
+ array_core_block4
x6 net46 net47 net48[9] net48[8] net48[7] net48[6] net48[5] net48[4] net48[3] net48[2] net48[1] net48[0] net49[9] net49[8]
+ net49[7] net49[6] net49[5] net49[4] net49[3] net49[2] net49[1] net49[0] net50[9] net50[8] net50[7] net50[6] net50[5] net50[4] net50[3]
+ net50[2] net50[1] net50[0] net51 net52 net53 net54[9] net54[8] net54[7] net54[6] net54[5] net54[4] net54[3] net54[2] net54[1] net54[0]
+ array_core_block5
x7 net55 net56 net57[4] net57[3] net57[2] net57[1] net57[0] net58[31] net58[30] net58[29] net58[28] net58[27] net58[26] net58[25]
+ net58[24] net58[23] net58[22] net58[21] net58[20] net58[19] net58[18] net58[17] net58[16] net58[15] net58[14] net58[13] net58[12] net58[11]
+ net58[10] net58[9] net58[8] net58[7] net58[6] net58[5] net58[4] net58[3] net58[2] net58[1] net58[0] array_row_decode
x8 net59 net60 net61[4] net61[3] net61[2] net61[1] net61[0] net62[31] net62[30] net62[29] net62[28] net62[27] net62[26] net62[25]
+ net62[24] net62[23] net62[22] net62[21] net62[20] net62[19] net62[18] net62[17] net62[16] net62[15] net62[14] net62[13] net62[12] net62[11]
+ net62[10] net62[9] net62[8] net62[7] net62[6] net62[5] net62[4] net62[3] net62[2] net62[1] net62[0] array_row_decode
.ends


* expanding   symbol:  array_core_block0.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block0.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block0.sch
.subckt array_core_block0 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_core_block1.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block1.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block1.sch
.subckt array_core_block1 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_core_block2.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block2.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block2.sch
.subckt array_core_block2 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_core_block3.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block3.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block3.sch
.subckt array_core_block3 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_core_block4.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block4.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block4.sch
.subckt array_core_block4 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_core_block5.sym # of pins=9
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block5.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_core_block5.sch
.subckt array_core_block5 vinj VGND vsrc[9] vsrc[8] vsrc[7] vsrc[6] vsrc[5] vsrc[4] vsrc[3] vsrc[2] vsrc[1] vsrc[0] row_en_6v0[9]
+ row_en_6v0[8] row_en_6v0[7] row_en_6v0[6] row_en_6v0[5] row_en_6v0[4] row_en_6v0[3] row_en_6v0[2] row_en_6v0[1] row_en_6v0[0] row_en_6v0_b[9]
+ row_en_6v0_b[8] row_en_6v0_b[7] row_en_6v0_b[6] row_en_6v0_b[5] row_en_6v0_b[4] row_en_6v0_b[3] row_en_6v0_b[2] row_en_6v0_b[1] row_en_6v0_b[0]
+ vtun vb vctrl vout[9] vout[8] vout[7] vout[6] vout[5] vout[4] vout[3] vout[2] vout[1] vout[0]
*.PININFO vtun:I vinj:I VGND:I vb:I row_en_6v0[9:0]:I row_en_6v0_b[9:0]:I vctrl:I vsrc[9:0]:I vout[9:0]:O
xc0[9] vb row_en_6v0[9] vinj vout[0] row_en_6v0_b[9] vtun vctrl vsrc[0] VGND net1[9] fgcell_amp
xc0[8] vb row_en_6v0[8] vinj vout[0] row_en_6v0_b[8] vtun vctrl vsrc[0] VGND net1[8] fgcell_amp
xc0[7] vb row_en_6v0[7] vinj vout[0] row_en_6v0_b[7] vtun vctrl vsrc[0] VGND net1[7] fgcell_amp
xc0[6] vb row_en_6v0[6] vinj vout[0] row_en_6v0_b[6] vtun vctrl vsrc[0] VGND net1[6] fgcell_amp
xc0[5] vb row_en_6v0[5] vinj vout[0] row_en_6v0_b[5] vtun vctrl vsrc[0] VGND net1[5] fgcell_amp
xc0[4] vb row_en_6v0[4] vinj vout[0] row_en_6v0_b[4] vtun vctrl vsrc[0] VGND net1[4] fgcell_amp
xc0[3] vb row_en_6v0[3] vinj vout[0] row_en_6v0_b[3] vtun vctrl vsrc[0] VGND net1[3] fgcell_amp
xc0[2] vb row_en_6v0[2] vinj vout[0] row_en_6v0_b[2] vtun vctrl vsrc[0] VGND net1[2] fgcell_amp
xc0[1] vb row_en_6v0[1] vinj vout[0] row_en_6v0_b[1] vtun vctrl vsrc[0] VGND net1[1] fgcell_amp
xc0[0] vb row_en_6v0[0] vinj vout[0] row_en_6v0_b[0] vtun vctrl vsrc[0] VGND net1[0] fgcell_amp
xc1[9] vb row_en_6v0[9] vinj vout[1] row_en_6v0_b[9] vtun vctrl vsrc[1] VGND net2[9] fgcell_amp
xc1[8] vb row_en_6v0[8] vinj vout[1] row_en_6v0_b[8] vtun vctrl vsrc[1] VGND net2[8] fgcell_amp
xc1[7] vb row_en_6v0[7] vinj vout[1] row_en_6v0_b[7] vtun vctrl vsrc[1] VGND net2[7] fgcell_amp
xc1[6] vb row_en_6v0[6] vinj vout[1] row_en_6v0_b[6] vtun vctrl vsrc[1] VGND net2[6] fgcell_amp
xc1[5] vb row_en_6v0[5] vinj vout[1] row_en_6v0_b[5] vtun vctrl vsrc[1] VGND net2[5] fgcell_amp
xc1[4] vb row_en_6v0[4] vinj vout[1] row_en_6v0_b[4] vtun vctrl vsrc[1] VGND net2[4] fgcell_amp
xc1[3] vb row_en_6v0[3] vinj vout[1] row_en_6v0_b[3] vtun vctrl vsrc[1] VGND net2[3] fgcell_amp
xc1[2] vb row_en_6v0[2] vinj vout[1] row_en_6v0_b[2] vtun vctrl vsrc[1] VGND net2[2] fgcell_amp
xc1[1] vb row_en_6v0[1] vinj vout[1] row_en_6v0_b[1] vtun vctrl vsrc[1] VGND net2[1] fgcell_amp
xc1[0] vb row_en_6v0[0] vinj vout[1] row_en_6v0_b[0] vtun vctrl vsrc[1] VGND net2[0] fgcell_amp
xc2[9] vb row_en_6v0[9] vinj vout[2] row_en_6v0_b[9] vtun vctrl vsrc[2] VGND net3[9] fgcell_amp
xc2[8] vb row_en_6v0[8] vinj vout[2] row_en_6v0_b[8] vtun vctrl vsrc[2] VGND net3[8] fgcell_amp
xc2[7] vb row_en_6v0[7] vinj vout[2] row_en_6v0_b[7] vtun vctrl vsrc[2] VGND net3[7] fgcell_amp
xc2[6] vb row_en_6v0[6] vinj vout[2] row_en_6v0_b[6] vtun vctrl vsrc[2] VGND net3[6] fgcell_amp
xc2[5] vb row_en_6v0[5] vinj vout[2] row_en_6v0_b[5] vtun vctrl vsrc[2] VGND net3[5] fgcell_amp
xc2[4] vb row_en_6v0[4] vinj vout[2] row_en_6v0_b[4] vtun vctrl vsrc[2] VGND net3[4] fgcell_amp
xc2[3] vb row_en_6v0[3] vinj vout[2] row_en_6v0_b[3] vtun vctrl vsrc[2] VGND net3[3] fgcell_amp
xc2[2] vb row_en_6v0[2] vinj vout[2] row_en_6v0_b[2] vtun vctrl vsrc[2] VGND net3[2] fgcell_amp
xc2[1] vb row_en_6v0[1] vinj vout[2] row_en_6v0_b[1] vtun vctrl vsrc[2] VGND net3[1] fgcell_amp
xc2[0] vb row_en_6v0[0] vinj vout[2] row_en_6v0_b[0] vtun vctrl vsrc[2] VGND net3[0] fgcell_amp
xc3[9] vb row_en_6v0[9] vinj vout[3] row_en_6v0_b[9] vtun vctrl vsrc[3] VGND net4[9] fgcell_amp
xc3[8] vb row_en_6v0[8] vinj vout[3] row_en_6v0_b[8] vtun vctrl vsrc[3] VGND net4[8] fgcell_amp
xc3[7] vb row_en_6v0[7] vinj vout[3] row_en_6v0_b[7] vtun vctrl vsrc[3] VGND net4[7] fgcell_amp
xc3[6] vb row_en_6v0[6] vinj vout[3] row_en_6v0_b[6] vtun vctrl vsrc[3] VGND net4[6] fgcell_amp
xc3[5] vb row_en_6v0[5] vinj vout[3] row_en_6v0_b[5] vtun vctrl vsrc[3] VGND net4[5] fgcell_amp
xc3[4] vb row_en_6v0[4] vinj vout[3] row_en_6v0_b[4] vtun vctrl vsrc[3] VGND net4[4] fgcell_amp
xc3[3] vb row_en_6v0[3] vinj vout[3] row_en_6v0_b[3] vtun vctrl vsrc[3] VGND net4[3] fgcell_amp
xc3[2] vb row_en_6v0[2] vinj vout[3] row_en_6v0_b[2] vtun vctrl vsrc[3] VGND net4[2] fgcell_amp
xc3[1] vb row_en_6v0[1] vinj vout[3] row_en_6v0_b[1] vtun vctrl vsrc[3] VGND net4[1] fgcell_amp
xc3[0] vb row_en_6v0[0] vinj vout[3] row_en_6v0_b[0] vtun vctrl vsrc[3] VGND net4[0] fgcell_amp
xc4[9] vb row_en_6v0[9] vinj vout[4] row_en_6v0_b[9] vtun vctrl vsrc[4] VGND net5[9] fgcell_amp
xc4[8] vb row_en_6v0[8] vinj vout[4] row_en_6v0_b[8] vtun vctrl vsrc[4] VGND net5[8] fgcell_amp
xc4[7] vb row_en_6v0[7] vinj vout[4] row_en_6v0_b[7] vtun vctrl vsrc[4] VGND net5[7] fgcell_amp
xc4[6] vb row_en_6v0[6] vinj vout[4] row_en_6v0_b[6] vtun vctrl vsrc[4] VGND net5[6] fgcell_amp
xc4[5] vb row_en_6v0[5] vinj vout[4] row_en_6v0_b[5] vtun vctrl vsrc[4] VGND net5[5] fgcell_amp
xc4[4] vb row_en_6v0[4] vinj vout[4] row_en_6v0_b[4] vtun vctrl vsrc[4] VGND net5[4] fgcell_amp
xc4[3] vb row_en_6v0[3] vinj vout[4] row_en_6v0_b[3] vtun vctrl vsrc[4] VGND net5[3] fgcell_amp
xc4[2] vb row_en_6v0[2] vinj vout[4] row_en_6v0_b[2] vtun vctrl vsrc[4] VGND net5[2] fgcell_amp
xc4[1] vb row_en_6v0[1] vinj vout[4] row_en_6v0_b[1] vtun vctrl vsrc[4] VGND net5[1] fgcell_amp
xc4[0] vb row_en_6v0[0] vinj vout[4] row_en_6v0_b[0] vtun vctrl vsrc[4] VGND net5[0] fgcell_amp
xc5[9] vb row_en_6v0[9] vinj vout[5] row_en_6v0_b[9] vtun vctrl vsrc[5] VGND net6[9] fgcell_amp
xc5[8] vb row_en_6v0[8] vinj vout[5] row_en_6v0_b[8] vtun vctrl vsrc[5] VGND net6[8] fgcell_amp
xc5[7] vb row_en_6v0[7] vinj vout[5] row_en_6v0_b[7] vtun vctrl vsrc[5] VGND net6[7] fgcell_amp
xc5[6] vb row_en_6v0[6] vinj vout[5] row_en_6v0_b[6] vtun vctrl vsrc[5] VGND net6[6] fgcell_amp
xc5[5] vb row_en_6v0[5] vinj vout[5] row_en_6v0_b[5] vtun vctrl vsrc[5] VGND net6[5] fgcell_amp
xc5[4] vb row_en_6v0[4] vinj vout[5] row_en_6v0_b[4] vtun vctrl vsrc[5] VGND net6[4] fgcell_amp
xc5[3] vb row_en_6v0[3] vinj vout[5] row_en_6v0_b[3] vtun vctrl vsrc[5] VGND net6[3] fgcell_amp
xc5[2] vb row_en_6v0[2] vinj vout[5] row_en_6v0_b[2] vtun vctrl vsrc[5] VGND net6[2] fgcell_amp
xc5[1] vb row_en_6v0[1] vinj vout[5] row_en_6v0_b[1] vtun vctrl vsrc[5] VGND net6[1] fgcell_amp
xc5[0] vb row_en_6v0[0] vinj vout[5] row_en_6v0_b[0] vtun vctrl vsrc[5] VGND net6[0] fgcell_amp
xc6[9] vb row_en_6v0[9] vinj vout[6] row_en_6v0_b[9] vtun vctrl vsrc[6] VGND net7[9] fgcell_amp
xc6[8] vb row_en_6v0[8] vinj vout[6] row_en_6v0_b[8] vtun vctrl vsrc[6] VGND net7[8] fgcell_amp
xc6[7] vb row_en_6v0[7] vinj vout[6] row_en_6v0_b[7] vtun vctrl vsrc[6] VGND net7[7] fgcell_amp
xc6[6] vb row_en_6v0[6] vinj vout[6] row_en_6v0_b[6] vtun vctrl vsrc[6] VGND net7[6] fgcell_amp
xc6[5] vb row_en_6v0[5] vinj vout[6] row_en_6v0_b[5] vtun vctrl vsrc[6] VGND net7[5] fgcell_amp
xc6[4] vb row_en_6v0[4] vinj vout[6] row_en_6v0_b[4] vtun vctrl vsrc[6] VGND net7[4] fgcell_amp
xc6[3] vb row_en_6v0[3] vinj vout[6] row_en_6v0_b[3] vtun vctrl vsrc[6] VGND net7[3] fgcell_amp
xc6[2] vb row_en_6v0[2] vinj vout[6] row_en_6v0_b[2] vtun vctrl vsrc[6] VGND net7[2] fgcell_amp
xc6[1] vb row_en_6v0[1] vinj vout[6] row_en_6v0_b[1] vtun vctrl vsrc[6] VGND net7[1] fgcell_amp
xc6[0] vb row_en_6v0[0] vinj vout[6] row_en_6v0_b[0] vtun vctrl vsrc[6] VGND net7[0] fgcell_amp
xc7[9] vb row_en_6v0[9] vinj vout[7] row_en_6v0_b[9] vtun vctrl vsrc[7] VGND net8[9] fgcell_amp
xc7[8] vb row_en_6v0[8] vinj vout[7] row_en_6v0_b[8] vtun vctrl vsrc[7] VGND net8[8] fgcell_amp
xc7[7] vb row_en_6v0[7] vinj vout[7] row_en_6v0_b[7] vtun vctrl vsrc[7] VGND net8[7] fgcell_amp
xc7[6] vb row_en_6v0[6] vinj vout[7] row_en_6v0_b[6] vtun vctrl vsrc[7] VGND net8[6] fgcell_amp
xc7[5] vb row_en_6v0[5] vinj vout[7] row_en_6v0_b[5] vtun vctrl vsrc[7] VGND net8[5] fgcell_amp
xc7[4] vb row_en_6v0[4] vinj vout[7] row_en_6v0_b[4] vtun vctrl vsrc[7] VGND net8[4] fgcell_amp
xc7[3] vb row_en_6v0[3] vinj vout[7] row_en_6v0_b[3] vtun vctrl vsrc[7] VGND net8[3] fgcell_amp
xc7[2] vb row_en_6v0[2] vinj vout[7] row_en_6v0_b[2] vtun vctrl vsrc[7] VGND net8[2] fgcell_amp
xc7[1] vb row_en_6v0[1] vinj vout[7] row_en_6v0_b[1] vtun vctrl vsrc[7] VGND net8[1] fgcell_amp
xc7[0] vb row_en_6v0[0] vinj vout[7] row_en_6v0_b[0] vtun vctrl vsrc[7] VGND net8[0] fgcell_amp
xc8[9] vb row_en_6v0[9] vinj vout[8] row_en_6v0_b[9] vtun vctrl vsrc[8] VGND net9[9] fgcell_amp
xc8[8] vb row_en_6v0[8] vinj vout[8] row_en_6v0_b[8] vtun vctrl vsrc[8] VGND net9[8] fgcell_amp
xc8[7] vb row_en_6v0[7] vinj vout[8] row_en_6v0_b[7] vtun vctrl vsrc[8] VGND net9[7] fgcell_amp
xc8[6] vb row_en_6v0[6] vinj vout[8] row_en_6v0_b[6] vtun vctrl vsrc[8] VGND net9[6] fgcell_amp
xc8[5] vb row_en_6v0[5] vinj vout[8] row_en_6v0_b[5] vtun vctrl vsrc[8] VGND net9[5] fgcell_amp
xc8[4] vb row_en_6v0[4] vinj vout[8] row_en_6v0_b[4] vtun vctrl vsrc[8] VGND net9[4] fgcell_amp
xc8[3] vb row_en_6v0[3] vinj vout[8] row_en_6v0_b[3] vtun vctrl vsrc[8] VGND net9[3] fgcell_amp
xc8[2] vb row_en_6v0[2] vinj vout[8] row_en_6v0_b[2] vtun vctrl vsrc[8] VGND net9[2] fgcell_amp
xc8[1] vb row_en_6v0[1] vinj vout[8] row_en_6v0_b[1] vtun vctrl vsrc[8] VGND net9[1] fgcell_amp
xc8[0] vb row_en_6v0[0] vinj vout[8] row_en_6v0_b[0] vtun vctrl vsrc[8] VGND net9[0] fgcell_amp
xc9[9] vb row_en_6v0[9] vinj vout[9] row_en_6v0_b[9] vtun vctrl vsrc[9] VGND net10[9] fgcell_amp
xc9[8] vb row_en_6v0[8] vinj vout[9] row_en_6v0_b[8] vtun vctrl vsrc[9] VGND net10[8] fgcell_amp
xc9[7] vb row_en_6v0[7] vinj vout[9] row_en_6v0_b[7] vtun vctrl vsrc[9] VGND net10[7] fgcell_amp
xc9[6] vb row_en_6v0[6] vinj vout[9] row_en_6v0_b[6] vtun vctrl vsrc[9] VGND net10[6] fgcell_amp
xc9[5] vb row_en_6v0[5] vinj vout[9] row_en_6v0_b[5] vtun vctrl vsrc[9] VGND net10[5] fgcell_amp
xc9[4] vb row_en_6v0[4] vinj vout[9] row_en_6v0_b[4] vtun vctrl vsrc[9] VGND net10[4] fgcell_amp
xc9[3] vb row_en_6v0[3] vinj vout[9] row_en_6v0_b[3] vtun vctrl vsrc[9] VGND net10[3] fgcell_amp
xc9[2] vb row_en_6v0[2] vinj vout[9] row_en_6v0_b[2] vtun vctrl vsrc[9] VGND net10[2] fgcell_amp
xc9[1] vb row_en_6v0[1] vinj vout[9] row_en_6v0_b[1] vtun vctrl vsrc[9] VGND net10[1] fgcell_amp
xc9[0] vb row_en_6v0[0] vinj vout[9] row_en_6v0_b[0] vtun vctrl vsrc[9] VGND net10[0] fgcell_amp
.ends


* expanding   symbol:  array_row_decode.sym # of pins=4
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_row_decode.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/array_row_decode.sch
.subckt array_row_decode VPWR VGND a[4] a[3] a[2] a[1] a[0] w[31] w[30] w[29] w[28] w[27] w[26] w[25] w[24] w[23] w[22] w[21]
+ w[20] w[19] w[18] w[17] w[16] w[15] w[14] w[13] w[12] w[11] w[10] w[9] w[8] w[7] w[6] w[5] w[4] w[3] w[2] w[1] w[0]
*.PININFO a[4:0]:I VPWR:I VGND:I w[31:0]:O
x1 a[4] VGND VGND VPWR VPWR net1 rowdec_not
x2 a[3] VGND VGND VPWR VPWR net2 rowdec_not
x3 a[2] VGND VGND VPWR VPWR net3 rowdec_not
x4 a[1] VGND VGND VPWR VPWR net4 rowdec_not
x5 a[0] VGND VGND VPWR VPWR net5 rowdec_not
x6 net5 net4 VGND VGND VPWR VPWR net6 rowdec_nand2
x7 a[0] net4 VGND VGND VPWR VPWR net8 rowdec_nand2
x8 net5 a[1] VGND VGND VPWR VPWR net9 rowdec_nand2
x9 a[0] a[1] VGND VGND VPWR VPWR net10 rowdec_nand2
x10 net3 net2 VGND VGND VPWR VPWR net7 rowdec_nand2
x11 a[2] net2 VGND VGND VPWR VPWR net11 rowdec_nand2
x12 net3 a[3] VGND VGND VPWR VPWR net12 rowdec_nand2
x13 a[2] a[3] VGND VGND VPWR VPWR net13 rowdec_nand2
x14 net6 net7 a[4] VGND VNB VPB VPWR w[0] rowdec_nor3
x15 net8 net7 a[4] VGND VNB VPB VPWR w[1] rowdec_nor3
x16 net9 net7 a[4] VGND VNB VPB VPWR w[2] rowdec_nor3
x17 net10 net7 a[4] VGND VNB VPB VPWR w[3] rowdec_nor3
x18 net6 net11 a[4] VGND VNB VPB VPWR w[4] rowdec_nor3
x19 net8 net11 a[4] VGND VNB VPB VPWR w[5] rowdec_nor3
x20 net9 net11 a[4] VGND VNB VPB VPWR w[6] rowdec_nor3
x21 net10 net11 a[4] VGND VNB VPB VPWR w[7] rowdec_nor3
x22 net6 net12 a[4] VGND VNB VPB VPWR w[8] rowdec_nor3
x23 net8 net12 a[4] VGND VNB VPB VPWR w[9] rowdec_nor3
x24 net9 net12 a[4] VGND VNB VPB VPWR w[10] rowdec_nor3
x25 net10 net12 a[4] VGND VNB VPB VPWR w[11] rowdec_nor3
x26 net6 net13 a[4] VGND VNB VPB VPWR w[12] rowdec_nor3
x27 net8 net13 a[4] VGND VNB VPB VPWR w[13] rowdec_nor3
x28 net9 net13 a[4] VGND VNB VPB VPWR w[14] rowdec_nor3
x29 net10 net13 a[4] VGND VNB VPB VPWR w[15] rowdec_nor3
x30 net6 net7 net1 VGND VNB VPB VPWR w[16] rowdec_nor3
x31 net8 net7 net1 VGND VNB VPB VPWR w[17] rowdec_nor3
x32 net9 net7 net1 VGND VNB VPB VPWR w[18] rowdec_nor3
x33 net10 net7 net1 VGND VNB VPB VPWR w[19] rowdec_nor3
x34 net6 net11 net1 VGND VNB VPB VPWR w[20] rowdec_nor3
x35 net8 net11 net1 VGND VNB VPB VPWR w[21] rowdec_nor3
x36 net9 net11 net1 VGND VNB VPB VPWR w[22] rowdec_nor3
x37 net10 net11 net1 VGND VNB VPB VPWR w[23] rowdec_nor3
x38 net6 net12 net1 VGND VNB VPB VPWR w[24] rowdec_nor3
x39 net8 net12 net1 VGND VNB VPB VPWR w[25] rowdec_nor3
x40 net9 net12 net1 VGND VNB VPB VPWR w[26] rowdec_nor3
x41 net10 net12 net1 VGND VNB VPB VPWR w[27] rowdec_nor3
x42 net6 net13 net1 VGND VNB VPB VPWR w[28] rowdec_nor3
x43 net8 net13 net1 VGND VNB VPB VPWR w[29] rowdec_nor3
x44 net9 net13 net1 VGND VNB VPB VPWR w[30] rowdec_nor3
x45 net10 net13 net1 VGND VNB VPB VPWR w[31] rowdec_nor3
.ends


* expanding   symbol:  fgcell_amp.sym # of pins=10
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/fgcell_amp.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/fgcell_amp.sch
.subckt fgcell_amp vb row_en_6v0 vinj vout row_en_6v0_b vtun vctrl vsrc VGND vfg
*.PININFO vinj:I row_en_6v0_b:I vtun:I vctrl:I vsrc:I vb:I VGND:I vout:O vfg:B row_en_6v0:I
x3 net1 vout row_en_6v0 row_en_6v0_b ideal_tg6v0
x1 vctrl vtun vinj row_en_6v0_b vsrc vfg VGND fgcell
x2 vinj vb net1 vfg net1 VGND diffamp_nmos
.ends


* expanding   symbol:  rowdec_not.sym # of pins=2
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_not.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_not.sch
.subckt rowdec_not A VGND VNB VPB VPWR Y
*.PININFO A:I Y:O
XM1 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  rowdec_nand2.sym # of pins=3
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_nand2.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_nand2.sch
.subckt rowdec_nand2 A B VGND VNB VPB VPWR Y
*.PININFO A:I Y:O B:I
XM1 Y A net1 VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net1 B VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  rowdec_nor3.sym # of pins=4
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_nor3.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/rowdec_nor3.sch
.subckt rowdec_nor3 A B C VGND VNB VPB VPWR Y
*.PININFO A:I Y:O B:I C:I
XM1 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 A VPWR VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 Y C VGND VNB sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net1 B net2 VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Y C net1 VPB sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  ideal_tg6v0.sym # of pins=4
** sym_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/ideal_tg6v0.sym
** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/ideal_tg6v0.sch
.subckt ideal_tg6v0 vin vout en en_b
*.PININFO vin:I en_b:I vout:O en:I
**** begin user architecture code


.model sw_vinj SW vt=3 vh=0.1 ron=14k roff=10gig
.model sw_1v8 SW vt={1.8/2}  vh=0.1 ron=10k roff=10gig


**** end user architecture code
S1 vin vout en en_b sw_vinj
.ends

.end
