magic
tech sky130A
timestamp 1717598570
<< pwell >>
rect 3300 19900 4441 21090
rect 15400 19900 16541 21090
<< psubdiff >>
rect 3300 21070 3312 21090
rect 4428 21070 4440 21090
rect 15400 21070 15412 21090
rect 16528 21070 16540 21090
<< psubdiffcont >>
rect 3312 21070 4428 21090
rect 15412 21070 16528 21090
<< locali >>
rect 3300 21070 3312 21090
rect 4428 21070 4440 21090
rect 15400 21070 15412 21090
rect 16528 21070 16540 21090
<< viali >>
rect 3312 21070 4428 21087
rect 15412 21072 16528 21089
<< metal1 >>
rect 3256 44021 3306 44024
rect 3256 43963 3259 44021
rect 3303 43963 3306 44021
rect 3256 41642 3306 43963
rect 16654 44021 16704 44024
rect 16654 43963 16657 44021
rect 16701 43963 16704 44021
rect 3256 41584 3259 41642
rect 3303 41584 3306 41642
rect 3256 41581 3306 41584
rect 3320 43931 3370 43934
rect 3320 43873 3323 43931
rect 3367 43873 3370 43931
rect 3320 41578 3370 43873
rect 16590 43931 16640 43934
rect 16590 43873 16593 43931
rect 16637 43873 16640 43931
rect 3320 41520 3323 41578
rect 3367 41520 3370 41578
rect 3320 41517 3370 41520
rect 3384 42521 3434 42524
rect 3384 42463 3387 42521
rect 3431 42463 3434 42521
rect 3384 41242 3434 42463
rect 16526 42521 16576 42524
rect 16526 42463 16529 42521
rect 16573 42463 16576 42521
rect 3384 41184 3387 41242
rect 3431 41184 3434 41242
rect 3384 41181 3434 41184
rect 3448 42431 3498 42434
rect 3448 42373 3451 42431
rect 3495 42373 3498 42431
rect 3448 41178 3498 42373
rect 16462 42431 16512 42434
rect 16462 42373 16465 42431
rect 16509 42373 16512 42431
rect 5087 41871 5173 41873
rect 5087 41793 5090 41871
rect 5170 41793 5173 41871
rect 14787 41871 14873 41873
rect 14787 41793 14790 41871
rect 14870 41793 14873 41871
rect 5090 41767 5170 41793
rect 3720 41725 5170 41767
rect 3677 41642 3727 41645
rect 3677 41598 3680 41642
rect 3724 41598 3727 41642
rect 3677 41595 3727 41598
rect 4989 41587 5047 41590
rect 3677 41578 3727 41581
rect 3677 41534 3680 41578
rect 3724 41534 3727 41578
rect 3677 41531 3727 41534
rect 4989 41535 4992 41587
rect 5044 41535 5047 41587
rect 4989 41532 5047 41535
rect 5031 41496 5063 41499
rect 3850 41447 3853 41473
rect 4257 41447 4260 41473
rect 3850 41444 4260 41447
rect 5031 41438 5034 41496
rect 5060 41438 5063 41496
rect 5031 41435 5063 41438
rect 5090 41367 5170 41725
rect 14790 41767 14870 41793
rect 14790 41725 16240 41767
rect 3673 41325 5170 41367
rect 3677 41242 3727 41245
rect 3677 41198 3680 41242
rect 3724 41198 3727 41242
rect 3677 41195 3727 41198
rect 4989 41187 5047 41190
rect 3448 41120 3451 41178
rect 3495 41120 3498 41178
rect 3677 41178 3727 41181
rect 3677 41134 3680 41178
rect 3724 41134 3727 41178
rect 3677 41131 3727 41134
rect 4989 41135 4992 41187
rect 5044 41135 5047 41187
rect 4989 41132 5047 41135
rect 3448 41117 3498 41120
rect 5031 41096 5063 41099
rect 3850 41047 3853 41073
rect 4257 41047 4260 41073
rect 3850 41044 4260 41047
rect 5031 41038 5034 41096
rect 5060 41038 5063 41096
rect 5031 41035 5063 41038
rect 3512 41021 3562 41024
rect 3512 40963 3515 41021
rect 3559 40963 3562 41021
rect 5090 41018 5170 41325
rect 14790 41367 14870 41725
rect 16233 41642 16283 41645
rect 16233 41598 16236 41642
rect 16280 41598 16283 41642
rect 16233 41595 16283 41598
rect 14913 41587 14971 41590
rect 14913 41535 14916 41587
rect 14968 41535 14971 41587
rect 14913 41532 14971 41535
rect 16233 41578 16283 41581
rect 16233 41534 16236 41578
rect 16280 41534 16283 41578
rect 16233 41531 16283 41534
rect 14897 41496 14929 41499
rect 14897 41438 14900 41496
rect 14926 41438 14929 41496
rect 15700 41447 15703 41473
rect 16107 41447 16110 41473
rect 15700 41442 16110 41447
rect 14897 41435 14929 41438
rect 14790 41325 16287 41367
rect 14790 41018 14870 41325
rect 16233 41242 16283 41245
rect 16233 41198 16236 41242
rect 16280 41198 16283 41242
rect 16233 41195 16283 41198
rect 14913 41187 14971 41190
rect 14913 41135 14916 41187
rect 14968 41135 14971 41187
rect 14913 41132 14971 41135
rect 16233 41178 16283 41181
rect 16233 41134 16236 41178
rect 16280 41134 16283 41178
rect 16233 41131 16283 41134
rect 16462 41178 16512 42373
rect 16526 41242 16576 42463
rect 16590 41578 16640 43873
rect 16654 41642 16704 43963
rect 16654 41584 16657 41642
rect 16701 41584 16704 41642
rect 16654 41581 16704 41584
rect 16590 41520 16593 41578
rect 16637 41520 16640 41578
rect 16590 41517 16640 41520
rect 16526 41184 16529 41242
rect 16573 41184 16576 41242
rect 16526 41181 16576 41184
rect 16462 41120 16465 41178
rect 16509 41120 16512 41178
rect 16462 41117 16512 41120
rect 14897 41096 14929 41099
rect 14897 41038 14900 41096
rect 14926 41038 14929 41096
rect 15700 41047 15703 41073
rect 16107 41047 16110 41073
rect 15700 41042 16110 41047
rect 14897 41035 14929 41038
rect 5090 40967 5141 41018
rect 3512 40842 3562 40963
rect 3673 40960 5141 40967
rect 5167 40960 5170 41018
rect 14790 40960 14793 41018
rect 14819 40967 14870 41018
rect 16398 41021 16448 41024
rect 14819 40960 16287 40967
rect 3512 40784 3515 40842
rect 3559 40784 3562 40842
rect 3512 40781 3562 40784
rect 3576 40931 3626 40934
rect 3576 40873 3579 40931
rect 3623 40873 3626 40931
rect 3673 40925 5170 40960
rect 3576 40778 3626 40873
rect 3677 40842 3727 40845
rect 3677 40798 3680 40842
rect 3724 40798 3727 40842
rect 3677 40795 3727 40798
rect 4989 40787 5047 40790
rect 3576 40720 3579 40778
rect 3623 40720 3626 40778
rect 3677 40778 3727 40781
rect 3677 40734 3680 40778
rect 3724 40734 3727 40778
rect 3677 40731 3727 40734
rect 4989 40735 4992 40787
rect 5044 40735 5047 40787
rect 4989 40732 5047 40735
rect 3576 40717 3626 40720
rect 5031 40696 5063 40699
rect 3850 40647 3853 40673
rect 4257 40647 4260 40673
rect 3850 40644 4260 40647
rect 5031 40638 5034 40696
rect 5060 40638 5063 40696
rect 5031 40635 5063 40638
rect 5090 40567 5170 40925
rect 14790 40925 16287 40960
rect 16398 40963 16401 41021
rect 16445 40963 16448 41021
rect 16334 40931 16384 40934
rect 3673 40525 5170 40567
rect 3576 40456 3626 40459
rect 3576 40398 3579 40456
rect 3623 40398 3626 40456
rect 3512 40392 3562 40395
rect 3512 40334 3515 40392
rect 3559 40334 3562 40392
rect 3448 40056 3498 40059
rect 3448 39998 3451 40056
rect 3495 39998 3498 40056
rect 3384 39992 3434 39995
rect 3384 39934 3387 39992
rect 3431 39934 3434 39992
rect 3320 39656 3370 39659
rect 3320 39598 3323 39656
rect 3367 39598 3370 39656
rect 3256 39592 3306 39595
rect 3256 39534 3259 39592
rect 3303 39534 3306 39592
rect 3192 39256 3242 39259
rect 3192 39198 3195 39256
rect 3239 39198 3242 39256
rect 3128 39192 3178 39195
rect 3128 39134 3131 39192
rect 3175 39134 3178 39192
rect 3064 38856 3114 38859
rect 3064 38798 3067 38856
rect 3111 38798 3114 38856
rect 3000 38792 3050 38795
rect 3000 38734 3003 38792
rect 3047 38734 3050 38792
rect 2936 38456 2986 38459
rect 2936 38398 2939 38456
rect 2983 38398 2986 38456
rect 2872 38392 2922 38395
rect 2872 38334 2875 38392
rect 2919 38334 2922 38392
rect 2808 38155 2858 38158
rect 2808 38097 2811 38155
rect 2855 38097 2858 38155
rect 2744 38091 2794 38094
rect 2744 38033 2747 38091
rect 2791 38033 2794 38091
rect 2680 37656 2730 37659
rect 2680 37598 2683 37656
rect 2727 37598 2730 37656
rect 2616 37592 2666 37595
rect 2616 37534 2619 37592
rect 2663 37534 2666 37592
rect 2552 37256 2602 37259
rect 2552 37198 2555 37256
rect 2599 37198 2602 37256
rect 2488 37192 2538 37195
rect 2488 37134 2491 37192
rect 2535 37134 2538 37192
rect 2424 36856 2474 36859
rect 2424 36798 2427 36856
rect 2471 36798 2474 36856
rect 2360 36792 2410 36795
rect 2360 36734 2363 36792
rect 2407 36734 2410 36792
rect 2296 36655 2346 36658
rect 2296 36597 2299 36655
rect 2343 36597 2346 36655
rect 2232 36591 2282 36594
rect 2232 36533 2235 36591
rect 2279 36533 2282 36591
rect 2168 36056 2218 36059
rect 2168 35998 2171 36056
rect 2215 35998 2218 36056
rect 2104 35992 2154 35995
rect 2104 35934 2107 35992
rect 2151 35934 2154 35992
rect 2040 35656 2090 35659
rect 2040 35598 2043 35656
rect 2087 35598 2090 35656
rect 1976 35592 2026 35595
rect 1976 35534 1979 35592
rect 2023 35534 2026 35592
rect 1912 35256 1962 35259
rect 1912 35198 1915 35256
rect 1959 35198 1962 35256
rect 1848 35192 1898 35195
rect 1848 35134 1851 35192
rect 1895 35134 1898 35192
rect 1784 34853 1834 34856
rect 1784 34795 1787 34853
rect 1831 34795 1834 34853
rect 1720 34789 1770 34792
rect 1720 34731 1723 34789
rect 1767 34731 1770 34789
rect 1656 34456 1706 34459
rect 1656 34398 1659 34456
rect 1703 34398 1706 34456
rect 1592 34392 1642 34395
rect 1592 34334 1595 34392
rect 1639 34334 1642 34392
rect 1528 34056 1578 34059
rect 1528 33998 1531 34056
rect 1575 33998 1578 34056
rect 1464 33992 1514 33995
rect 1464 33934 1467 33992
rect 1511 33934 1514 33992
rect 1400 33656 1450 33659
rect 1400 33598 1403 33656
rect 1447 33598 1450 33656
rect 1336 33592 1386 33595
rect 1336 33534 1339 33592
rect 1383 33534 1386 33592
rect 1272 33256 1322 33259
rect 1272 33198 1275 33256
rect 1319 33198 1322 33256
rect 1208 33192 1258 33195
rect 1208 33134 1211 33192
rect 1255 33134 1258 33192
rect 1144 32856 1194 32859
rect 1144 32798 1147 32856
rect 1191 32798 1194 32856
rect 1080 32792 1130 32795
rect 1080 32734 1083 32792
rect 1127 32734 1130 32792
rect 1016 32456 1066 32459
rect 1016 32398 1019 32456
rect 1063 32398 1066 32456
rect 952 32392 1002 32395
rect 952 32334 955 32392
rect 999 32334 1002 32392
rect 888 32149 938 32152
rect 888 32091 891 32149
rect 935 32091 938 32149
rect 824 32085 874 32088
rect 824 32027 827 32085
rect 871 32027 874 32085
rect 760 31656 810 31659
rect 760 31598 763 31656
rect 807 31598 810 31656
rect 696 31592 746 31595
rect 696 31534 699 31592
rect 743 31534 746 31592
rect 632 31256 682 31259
rect 632 31198 635 31256
rect 679 31198 682 31256
rect 568 31192 618 31195
rect 568 31134 571 31192
rect 615 31134 618 31192
rect 504 30856 554 30859
rect 504 30798 507 30856
rect 551 30798 554 30856
rect 440 30792 490 30795
rect 440 30734 443 30792
rect 487 30734 490 30792
rect 376 30655 426 30658
rect 376 30597 379 30655
rect 423 30597 426 30655
rect 312 30591 362 30594
rect 312 30533 315 30591
rect 359 30533 362 30591
rect 248 30056 298 30059
rect 248 29998 251 30056
rect 295 29998 298 30056
rect 184 29992 234 29995
rect 184 29934 187 29992
rect 231 29934 234 29992
rect 184 417 234 29934
rect 248 507 298 29998
rect 312 1917 362 30533
rect 376 2007 426 30597
rect 440 3417 490 30734
rect 504 3507 554 30798
rect 568 4917 618 31134
rect 632 5007 682 31198
rect 696 6417 746 31534
rect 760 6507 810 31598
rect 824 7917 874 32027
rect 888 8007 938 32091
rect 952 9417 1002 32334
rect 1016 9507 1066 32398
rect 1080 10917 1130 32734
rect 1144 11007 1194 32798
rect 1208 12417 1258 33134
rect 1272 12507 1322 33198
rect 1336 13917 1386 33534
rect 1400 14007 1450 33598
rect 1464 15417 1514 33934
rect 1528 15507 1578 33998
rect 1592 16917 1642 34334
rect 1656 17007 1706 34398
rect 1720 18417 1770 34731
rect 1784 18507 1834 34795
rect 1848 19917 1898 35134
rect 1912 20007 1962 35198
rect 1976 21417 2026 35534
rect 2040 21507 2090 35598
rect 2104 22917 2154 35934
rect 2168 23007 2218 35998
rect 2232 24417 2282 36533
rect 2296 24507 2346 36597
rect 2360 25917 2410 36734
rect 2424 26007 2474 36798
rect 2488 27417 2538 37134
rect 2552 27507 2602 37198
rect 2616 28917 2666 37534
rect 2680 29007 2730 37598
rect 2744 30417 2794 38033
rect 2808 30507 2858 38097
rect 2872 31917 2922 38334
rect 2936 32007 2986 38398
rect 3000 33417 3050 38734
rect 3064 33507 3114 38798
rect 3128 34917 3178 39134
rect 3192 35007 3242 39198
rect 3256 36417 3306 39534
rect 3320 36507 3370 39598
rect 3384 37917 3434 39934
rect 3448 38007 3498 39998
rect 3512 39417 3562 40334
rect 3576 39507 3626 40398
rect 3677 40442 3727 40445
rect 3677 40398 3680 40442
rect 3724 40398 3727 40442
rect 3677 40395 3727 40398
rect 4989 40387 5047 40390
rect 3677 40378 3727 40381
rect 3677 40334 3680 40378
rect 3724 40334 3727 40378
rect 3677 40331 3727 40334
rect 4989 40335 4992 40387
rect 5044 40335 5047 40387
rect 4989 40332 5047 40335
rect 5031 40296 5063 40299
rect 3850 40247 3853 40273
rect 4257 40247 4260 40273
rect 3850 40244 4260 40247
rect 5031 40238 5034 40296
rect 5060 40238 5063 40296
rect 5031 40235 5063 40238
rect 5090 40218 5170 40525
rect 14790 40567 14870 40925
rect 16334 40873 16337 40931
rect 16381 40873 16384 40931
rect 16233 40842 16283 40845
rect 16233 40798 16236 40842
rect 16280 40798 16283 40842
rect 16233 40795 16283 40798
rect 14913 40787 14971 40790
rect 14913 40735 14916 40787
rect 14968 40735 14971 40787
rect 14913 40732 14971 40735
rect 16233 40778 16283 40781
rect 16233 40734 16236 40778
rect 16280 40734 16283 40778
rect 16233 40731 16283 40734
rect 16334 40778 16384 40873
rect 16398 40842 16448 40963
rect 16398 40784 16401 40842
rect 16445 40784 16448 40842
rect 16398 40781 16448 40784
rect 16334 40720 16337 40778
rect 16381 40720 16384 40778
rect 16334 40717 16384 40720
rect 14897 40696 14929 40699
rect 14897 40638 14900 40696
rect 14926 40638 14929 40696
rect 15700 40647 15703 40673
rect 16107 40647 16110 40673
rect 15700 40642 16110 40647
rect 14897 40635 14929 40638
rect 14790 40525 16287 40567
rect 14790 40218 14870 40525
rect 16334 40456 16384 40459
rect 16233 40442 16283 40445
rect 16233 40398 16236 40442
rect 16280 40398 16283 40442
rect 16233 40395 16283 40398
rect 16334 40398 16337 40456
rect 16381 40398 16384 40456
rect 14913 40387 14971 40390
rect 14913 40335 14916 40387
rect 14968 40335 14971 40387
rect 14913 40332 14971 40335
rect 16233 40378 16283 40381
rect 16233 40334 16236 40378
rect 16280 40334 16283 40378
rect 16233 40331 16283 40334
rect 14897 40296 14929 40299
rect 14897 40238 14900 40296
rect 14926 40238 14929 40296
rect 15700 40247 15703 40273
rect 16107 40247 16110 40273
rect 15700 40242 16110 40247
rect 14897 40235 14929 40238
rect 5090 40167 5141 40218
rect 3673 40160 5141 40167
rect 5167 40160 5170 40218
rect 14790 40160 14793 40218
rect 14819 40167 14870 40218
rect 14819 40160 16287 40167
rect 3673 40125 5170 40160
rect 3677 40042 3727 40045
rect 3677 39998 3680 40042
rect 3724 39998 3727 40042
rect 3677 39995 3727 39998
rect 4989 39987 5047 39990
rect 3677 39978 3727 39981
rect 3677 39934 3680 39978
rect 3724 39934 3727 39978
rect 3677 39931 3727 39934
rect 4989 39935 4992 39987
rect 5044 39935 5047 39987
rect 4989 39932 5047 39935
rect 5031 39896 5063 39899
rect 3850 39847 3853 39873
rect 4257 39847 4260 39873
rect 3850 39844 4260 39847
rect 5031 39838 5034 39896
rect 5060 39838 5063 39896
rect 5031 39835 5063 39838
rect 5090 39767 5170 40125
rect 14790 40125 16287 40160
rect 3673 39725 5170 39767
rect 3677 39642 3727 39645
rect 3677 39598 3680 39642
rect 3724 39598 3727 39642
rect 3677 39595 3727 39598
rect 4989 39587 5047 39590
rect 3677 39578 3727 39581
rect 3677 39534 3680 39578
rect 3724 39534 3727 39578
rect 3677 39531 3727 39534
rect 4989 39535 4992 39587
rect 5044 39535 5047 39587
rect 4989 39532 5047 39535
rect 3576 39449 3579 39507
rect 3623 39449 3626 39507
rect 5031 39496 5063 39499
rect 3576 39446 3626 39449
rect 3850 39447 3853 39473
rect 4257 39447 4260 39473
rect 3850 39444 4260 39447
rect 5031 39438 5034 39496
rect 5060 39438 5063 39496
rect 5031 39435 5063 39438
rect 3512 39359 3515 39417
rect 3559 39359 3562 39417
rect 5090 39418 5170 39725
rect 14790 39767 14870 40125
rect 16233 40042 16283 40045
rect 16233 39998 16236 40042
rect 16280 39998 16283 40042
rect 16233 39995 16283 39998
rect 14913 39987 14971 39990
rect 14913 39935 14916 39987
rect 14968 39935 14971 39987
rect 14913 39932 14971 39935
rect 16233 39978 16283 39981
rect 16233 39934 16236 39978
rect 16280 39934 16283 39978
rect 16233 39931 16283 39934
rect 14897 39896 14929 39899
rect 14897 39838 14900 39896
rect 14926 39838 14929 39896
rect 15700 39847 15703 39873
rect 16107 39847 16110 39873
rect 15700 39842 16110 39847
rect 14897 39835 14929 39838
rect 14790 39725 16287 39767
rect 14790 39418 14870 39725
rect 16233 39642 16283 39645
rect 16233 39598 16236 39642
rect 16280 39598 16283 39642
rect 16233 39595 16283 39598
rect 14913 39587 14971 39590
rect 14913 39535 14916 39587
rect 14968 39535 14971 39587
rect 14913 39532 14971 39535
rect 16233 39578 16283 39581
rect 16233 39534 16236 39578
rect 16280 39534 16283 39578
rect 16233 39531 16283 39534
rect 16334 39507 16384 40398
rect 14897 39496 14929 39499
rect 14897 39438 14900 39496
rect 14926 39438 14929 39496
rect 15700 39447 15703 39473
rect 16107 39447 16110 39473
rect 15700 39442 16110 39447
rect 16334 39449 16337 39507
rect 16381 39449 16384 39507
rect 16334 39446 16384 39449
rect 16398 40392 16448 40395
rect 16398 40334 16401 40392
rect 16445 40334 16448 40392
rect 14897 39435 14929 39438
rect 5090 39367 5141 39418
rect 3512 39356 3562 39359
rect 3673 39360 5141 39367
rect 5167 39360 5170 39418
rect 14790 39360 14793 39418
rect 14819 39367 14870 39418
rect 16398 39417 16448 40334
rect 14819 39360 16287 39367
rect 3673 39325 5170 39360
rect 3677 39242 3727 39245
rect 3677 39198 3680 39242
rect 3724 39198 3727 39242
rect 3677 39195 3727 39198
rect 4989 39187 5047 39190
rect 3677 39178 3727 39181
rect 3677 39134 3680 39178
rect 3724 39134 3727 39178
rect 3677 39131 3727 39134
rect 4989 39135 4992 39187
rect 5044 39135 5047 39187
rect 4989 39132 5047 39135
rect 5031 39096 5063 39099
rect 3850 39047 3853 39073
rect 4257 39047 4260 39073
rect 3850 39044 4260 39047
rect 5031 39038 5034 39096
rect 5060 39038 5063 39096
rect 5031 39035 5063 39038
rect 5090 38967 5170 39325
rect 14790 39325 16287 39360
rect 16398 39359 16401 39417
rect 16445 39359 16448 39417
rect 16398 39356 16448 39359
rect 16462 40056 16512 40059
rect 16462 39998 16465 40056
rect 16509 39998 16512 40056
rect 3673 38925 5170 38967
rect 3677 38842 3727 38845
rect 3677 38798 3680 38842
rect 3724 38798 3727 38842
rect 3677 38795 3727 38798
rect 4989 38787 5047 38790
rect 3677 38778 3727 38781
rect 3677 38734 3680 38778
rect 3724 38734 3727 38778
rect 3677 38731 3727 38734
rect 4989 38735 4992 38787
rect 5044 38735 5047 38787
rect 4989 38732 5047 38735
rect 5031 38696 5063 38699
rect 3850 38647 3853 38673
rect 4257 38647 4260 38673
rect 3850 38644 4260 38647
rect 5031 38638 5034 38696
rect 5060 38638 5063 38696
rect 5031 38635 5063 38638
rect 5090 38618 5170 38925
rect 14790 38967 14870 39325
rect 16233 39242 16283 39245
rect 16233 39198 16236 39242
rect 16280 39198 16283 39242
rect 16233 39195 16283 39198
rect 14913 39187 14971 39190
rect 14913 39135 14916 39187
rect 14968 39135 14971 39187
rect 14913 39132 14971 39135
rect 16233 39178 16283 39181
rect 16233 39134 16236 39178
rect 16280 39134 16283 39178
rect 16233 39131 16283 39134
rect 14897 39096 14929 39099
rect 14897 39038 14900 39096
rect 14926 39038 14929 39096
rect 15700 39047 15703 39073
rect 16107 39047 16110 39073
rect 15700 39042 16110 39047
rect 14897 39035 14929 39038
rect 14790 38925 16287 38967
rect 14790 38618 14870 38925
rect 16233 38842 16283 38845
rect 16233 38798 16236 38842
rect 16280 38798 16283 38842
rect 16233 38795 16283 38798
rect 14913 38787 14971 38790
rect 14913 38735 14916 38787
rect 14968 38735 14971 38787
rect 14913 38732 14971 38735
rect 16233 38778 16283 38781
rect 16233 38734 16236 38778
rect 16280 38734 16283 38778
rect 16233 38731 16283 38734
rect 14897 38696 14929 38699
rect 14897 38638 14900 38696
rect 14926 38638 14929 38696
rect 15700 38647 15703 38673
rect 16107 38647 16110 38673
rect 15700 38642 16110 38647
rect 14897 38635 14929 38638
rect 5090 38567 5141 38618
rect 3673 38560 5141 38567
rect 5167 38560 5170 38618
rect 14790 38560 14793 38618
rect 14819 38567 14870 38618
rect 14819 38560 16287 38567
rect 3673 38525 5170 38560
rect 3677 38442 3727 38445
rect 3677 38398 3680 38442
rect 3724 38398 3727 38442
rect 3677 38395 3727 38398
rect 4989 38387 5047 38390
rect 3677 38378 3727 38381
rect 3677 38334 3680 38378
rect 3724 38334 3727 38378
rect 3677 38331 3727 38334
rect 4989 38335 4992 38387
rect 5044 38335 5047 38387
rect 4989 38332 5047 38335
rect 5031 38296 5063 38299
rect 3850 38247 3853 38273
rect 4257 38247 4260 38273
rect 3850 38244 4260 38247
rect 5031 38238 5034 38296
rect 5060 38238 5063 38296
rect 5031 38235 5063 38238
rect 5090 38167 5170 38525
rect 14790 38525 16287 38560
rect 3673 38125 5170 38167
rect 3448 37949 3451 38007
rect 3495 37949 3498 38007
rect 3677 38042 3727 38045
rect 3677 37998 3680 38042
rect 3724 37998 3727 38042
rect 3677 37995 3727 37998
rect 4989 37987 5047 37990
rect 3448 37946 3498 37949
rect 3677 37978 3727 37981
rect 3677 37934 3680 37978
rect 3724 37934 3727 37978
rect 3677 37931 3727 37934
rect 4989 37935 4992 37987
rect 5044 37935 5047 37987
rect 4989 37932 5047 37935
rect 3384 37859 3387 37917
rect 3431 37859 3434 37917
rect 5031 37896 5063 37899
rect 3384 37856 3434 37859
rect 3850 37847 3853 37873
rect 4257 37847 4260 37873
rect 3850 37844 4260 37847
rect 5031 37838 5034 37896
rect 5060 37838 5063 37896
rect 5031 37835 5063 37838
rect 5090 37818 5170 38125
rect 14790 38167 14870 38525
rect 16233 38442 16283 38445
rect 16233 38398 16236 38442
rect 16280 38398 16283 38442
rect 16233 38395 16283 38398
rect 14913 38387 14971 38390
rect 14913 38335 14916 38387
rect 14968 38335 14971 38387
rect 14913 38332 14971 38335
rect 16233 38378 16283 38381
rect 16233 38334 16236 38378
rect 16280 38334 16283 38378
rect 16233 38331 16283 38334
rect 14897 38296 14929 38299
rect 14897 38238 14900 38296
rect 14926 38238 14929 38296
rect 15700 38247 15703 38273
rect 16107 38247 16110 38273
rect 15700 38242 16110 38247
rect 14897 38235 14929 38238
rect 14790 38125 16287 38167
rect 14790 37818 14870 38125
rect 16233 38042 16283 38045
rect 16233 37998 16236 38042
rect 16280 37998 16283 38042
rect 16233 37995 16283 37998
rect 16462 38007 16512 39998
rect 14913 37987 14971 37990
rect 14913 37935 14916 37987
rect 14968 37935 14971 37987
rect 14913 37932 14971 37935
rect 16233 37978 16283 37981
rect 16233 37934 16236 37978
rect 16280 37934 16283 37978
rect 16462 37949 16465 38007
rect 16509 37949 16512 38007
rect 16462 37946 16512 37949
rect 16526 39992 16576 39995
rect 16526 39934 16529 39992
rect 16573 39934 16576 39992
rect 16233 37931 16283 37934
rect 16526 37917 16576 39934
rect 14897 37896 14929 37899
rect 14897 37838 14900 37896
rect 14926 37838 14929 37896
rect 15700 37847 15703 37873
rect 16107 37847 16110 37873
rect 16526 37859 16529 37917
rect 16573 37859 16576 37917
rect 16526 37856 16576 37859
rect 16590 39656 16640 39659
rect 16590 39598 16593 39656
rect 16637 39598 16640 39656
rect 15700 37842 16110 37847
rect 14897 37835 14929 37838
rect 5090 37767 5141 37818
rect 3673 37760 5141 37767
rect 5167 37760 5170 37818
rect 14790 37760 14793 37818
rect 14819 37767 14870 37818
rect 14819 37760 16287 37767
rect 3673 37725 5170 37760
rect 3677 37642 3727 37645
rect 3677 37598 3680 37642
rect 3724 37598 3727 37642
rect 3677 37595 3727 37598
rect 4989 37587 5047 37590
rect 3677 37578 3727 37581
rect 3677 37534 3680 37578
rect 3724 37534 3727 37578
rect 3677 37531 3727 37534
rect 4989 37535 4992 37587
rect 5044 37535 5047 37587
rect 4989 37532 5047 37535
rect 5031 37496 5063 37499
rect 3850 37447 3853 37473
rect 4257 37447 4260 37473
rect 3850 37444 4260 37447
rect 5031 37438 5034 37496
rect 5060 37438 5063 37496
rect 5031 37435 5063 37438
rect 5090 37367 5170 37725
rect 14790 37725 16287 37760
rect 3673 37325 5170 37367
rect 3677 37242 3727 37245
rect 3677 37198 3680 37242
rect 3724 37198 3727 37242
rect 3677 37195 3727 37198
rect 4989 37187 5047 37190
rect 3677 37178 3727 37181
rect 3677 37134 3680 37178
rect 3724 37134 3727 37178
rect 3677 37131 3727 37134
rect 4989 37135 4992 37187
rect 5044 37135 5047 37187
rect 4989 37132 5047 37135
rect 5031 37096 5063 37099
rect 3850 37047 3853 37073
rect 4257 37047 4260 37073
rect 3850 37044 4260 37047
rect 5031 37038 5034 37096
rect 5060 37038 5063 37096
rect 5031 37035 5063 37038
rect 5090 37018 5170 37325
rect 14790 37367 14870 37725
rect 16233 37642 16283 37645
rect 16233 37598 16236 37642
rect 16280 37598 16283 37642
rect 16233 37595 16283 37598
rect 14913 37587 14971 37590
rect 14913 37535 14916 37587
rect 14968 37535 14971 37587
rect 14913 37532 14971 37535
rect 16233 37578 16283 37581
rect 16233 37534 16236 37578
rect 16280 37534 16283 37578
rect 16233 37531 16283 37534
rect 14897 37496 14929 37499
rect 14897 37438 14900 37496
rect 14926 37438 14929 37496
rect 15700 37447 15703 37473
rect 16107 37447 16110 37473
rect 15700 37442 16110 37447
rect 14897 37435 14929 37438
rect 14790 37325 16287 37367
rect 14790 37018 14870 37325
rect 16233 37242 16283 37245
rect 16233 37198 16236 37242
rect 16280 37198 16283 37242
rect 16233 37195 16283 37198
rect 14913 37187 14971 37190
rect 14913 37135 14916 37187
rect 14968 37135 14971 37187
rect 14913 37132 14971 37135
rect 16233 37178 16283 37181
rect 16233 37134 16236 37178
rect 16280 37134 16283 37178
rect 16233 37131 16283 37134
rect 14897 37096 14929 37099
rect 14897 37038 14900 37096
rect 14926 37038 14929 37096
rect 15700 37047 15703 37073
rect 16107 37047 16110 37073
rect 15700 37042 16110 37047
rect 14897 37035 14929 37038
rect 5090 36967 5141 37018
rect 3673 36960 5141 36967
rect 5167 36960 5170 37018
rect 14790 36960 14793 37018
rect 14819 36967 14870 37018
rect 14819 36960 16287 36967
rect 3673 36925 5170 36960
rect 3677 36842 3727 36845
rect 3677 36798 3680 36842
rect 3724 36798 3727 36842
rect 3677 36795 3727 36798
rect 4989 36787 5047 36790
rect 3677 36778 3727 36781
rect 3677 36734 3680 36778
rect 3724 36734 3727 36778
rect 3677 36731 3727 36734
rect 4989 36735 4992 36787
rect 5044 36735 5047 36787
rect 4989 36732 5047 36735
rect 5031 36696 5063 36699
rect 3850 36647 3853 36673
rect 4257 36647 4260 36673
rect 3850 36644 4260 36647
rect 5031 36638 5034 36696
rect 5060 36638 5063 36696
rect 5031 36635 5063 36638
rect 5090 36567 5170 36925
rect 14790 36925 16287 36960
rect 3673 36525 5170 36567
rect 3320 36449 3323 36507
rect 3367 36449 3370 36507
rect 3320 36446 3370 36449
rect 3256 36359 3259 36417
rect 3303 36359 3306 36417
rect 3677 36442 3727 36445
rect 3677 36398 3680 36442
rect 3724 36398 3727 36442
rect 3677 36395 3727 36398
rect 4989 36387 5047 36390
rect 3256 36356 3306 36359
rect 3677 36378 3727 36381
rect 3677 36334 3680 36378
rect 3724 36334 3727 36378
rect 3677 36331 3727 36334
rect 4989 36335 4992 36387
rect 5044 36335 5047 36387
rect 4989 36332 5047 36335
rect 5031 36296 5063 36299
rect 3850 36247 3853 36273
rect 4257 36247 4260 36273
rect 3850 36244 4260 36247
rect 5031 36238 5034 36296
rect 5060 36238 5063 36296
rect 5031 36235 5063 36238
rect 5090 36218 5170 36525
rect 14790 36567 14870 36925
rect 16233 36842 16283 36845
rect 16233 36798 16236 36842
rect 16280 36798 16283 36842
rect 16233 36795 16283 36798
rect 14913 36787 14971 36790
rect 14913 36735 14916 36787
rect 14968 36735 14971 36787
rect 14913 36732 14971 36735
rect 16233 36778 16283 36781
rect 16233 36734 16236 36778
rect 16280 36734 16283 36778
rect 16233 36731 16283 36734
rect 14897 36696 14929 36699
rect 14897 36638 14900 36696
rect 14926 36638 14929 36696
rect 15700 36647 15703 36673
rect 16107 36647 16110 36673
rect 15700 36642 16110 36647
rect 14897 36635 14929 36638
rect 14790 36525 16287 36567
rect 14790 36218 14870 36525
rect 16590 36507 16640 39598
rect 16590 36449 16593 36507
rect 16637 36449 16640 36507
rect 16590 36446 16640 36449
rect 16654 39592 16704 39595
rect 16654 39534 16657 39592
rect 16701 39534 16704 39592
rect 16233 36442 16283 36445
rect 16233 36398 16236 36442
rect 16280 36398 16283 36442
rect 16233 36395 16283 36398
rect 16654 36417 16704 39534
rect 14913 36387 14971 36390
rect 14913 36335 14916 36387
rect 14968 36335 14971 36387
rect 14913 36332 14971 36335
rect 16233 36378 16283 36381
rect 16233 36334 16236 36378
rect 16280 36334 16283 36378
rect 16654 36359 16657 36417
rect 16701 36359 16704 36417
rect 16654 36356 16704 36359
rect 16718 39256 16768 39259
rect 16718 39198 16721 39256
rect 16765 39198 16768 39256
rect 16233 36331 16283 36334
rect 14897 36296 14929 36299
rect 14897 36238 14900 36296
rect 14926 36238 14929 36296
rect 15700 36247 15703 36273
rect 16107 36247 16110 36273
rect 15700 36242 16110 36247
rect 14897 36235 14929 36238
rect 5090 36167 5141 36218
rect 3673 36160 5141 36167
rect 5167 36160 5170 36218
rect 14790 36160 14793 36218
rect 14819 36167 14870 36218
rect 14819 36160 16287 36167
rect 3673 36125 5170 36160
rect 3677 36042 3727 36045
rect 3677 35998 3680 36042
rect 3724 35998 3727 36042
rect 3677 35995 3727 35998
rect 4989 35987 5047 35990
rect 3677 35978 3727 35981
rect 3677 35934 3680 35978
rect 3724 35934 3727 35978
rect 3677 35931 3727 35934
rect 4989 35935 4992 35987
rect 5044 35935 5047 35987
rect 4989 35932 5047 35935
rect 5031 35896 5063 35899
rect 3850 35847 3853 35873
rect 4257 35847 4260 35873
rect 3850 35844 4260 35847
rect 5031 35838 5034 35896
rect 5060 35838 5063 35896
rect 5031 35835 5063 35838
rect 5090 35767 5170 36125
rect 14790 36125 16287 36160
rect 3673 35725 5170 35767
rect 3677 35642 3727 35645
rect 3677 35598 3680 35642
rect 3724 35598 3727 35642
rect 3677 35595 3727 35598
rect 4989 35587 5047 35590
rect 3677 35578 3727 35581
rect 3677 35534 3680 35578
rect 3724 35534 3727 35578
rect 3677 35531 3727 35534
rect 4989 35535 4992 35587
rect 5044 35535 5047 35587
rect 4989 35532 5047 35535
rect 5031 35496 5063 35499
rect 3850 35447 3853 35473
rect 4257 35447 4260 35473
rect 3850 35444 4260 35447
rect 5031 35438 5034 35496
rect 5060 35438 5063 35496
rect 5031 35435 5063 35438
rect 5090 35418 5170 35725
rect 14790 35767 14870 36125
rect 16233 36042 16283 36045
rect 16233 35998 16236 36042
rect 16280 35998 16283 36042
rect 16233 35995 16283 35998
rect 14913 35987 14971 35990
rect 14913 35935 14916 35987
rect 14968 35935 14971 35987
rect 14913 35932 14971 35935
rect 16233 35978 16283 35981
rect 16233 35934 16236 35978
rect 16280 35934 16283 35978
rect 16233 35931 16283 35934
rect 14897 35896 14929 35899
rect 14897 35838 14900 35896
rect 14926 35838 14929 35896
rect 15700 35847 15703 35873
rect 16107 35847 16110 35873
rect 15700 35842 16110 35847
rect 14897 35835 14929 35838
rect 14790 35725 16287 35767
rect 14790 35418 14870 35725
rect 16233 35642 16283 35645
rect 16233 35598 16236 35642
rect 16280 35598 16283 35642
rect 16233 35595 16283 35598
rect 14913 35587 14971 35590
rect 14913 35535 14916 35587
rect 14968 35535 14971 35587
rect 14913 35532 14971 35535
rect 16233 35578 16283 35581
rect 16233 35534 16236 35578
rect 16280 35534 16283 35578
rect 16233 35531 16283 35534
rect 14897 35496 14929 35499
rect 14897 35438 14900 35496
rect 14926 35438 14929 35496
rect 15700 35447 15703 35473
rect 16107 35447 16110 35473
rect 15700 35442 16110 35447
rect 14897 35435 14929 35438
rect 5090 35367 5141 35418
rect 3673 35360 5141 35367
rect 5167 35360 5170 35418
rect 14790 35360 14793 35418
rect 14819 35367 14870 35418
rect 14819 35360 16287 35367
rect 3673 35325 5170 35360
rect 3677 35242 3727 35245
rect 3677 35198 3680 35242
rect 3724 35198 3727 35242
rect 3677 35195 3727 35198
rect 4989 35187 5047 35190
rect 3677 35178 3727 35181
rect 3677 35134 3680 35178
rect 3724 35134 3727 35178
rect 3677 35131 3727 35134
rect 4989 35135 4992 35187
rect 5044 35135 5047 35187
rect 4989 35132 5047 35135
rect 5031 35096 5063 35099
rect 3850 35047 3853 35073
rect 4257 35047 4260 35073
rect 3850 35044 4260 35047
rect 5031 35038 5034 35096
rect 5060 35038 5063 35096
rect 5031 35035 5063 35038
rect 3192 34949 3195 35007
rect 3239 34949 3242 35007
rect 5090 34967 5170 35325
rect 14790 35325 16287 35360
rect 3192 34946 3242 34949
rect 3673 34925 5170 34967
rect 3128 34859 3131 34917
rect 3175 34859 3178 34917
rect 3128 34856 3178 34859
rect 3677 34842 3727 34845
rect 3677 34798 3680 34842
rect 3724 34798 3727 34842
rect 3677 34795 3727 34798
rect 4989 34787 5047 34790
rect 3677 34778 3727 34781
rect 3677 34734 3680 34778
rect 3724 34734 3727 34778
rect 3677 34731 3727 34734
rect 4989 34735 4992 34787
rect 5044 34735 5047 34787
rect 4989 34732 5047 34735
rect 5031 34696 5063 34699
rect 3850 34647 3853 34673
rect 4257 34647 4260 34673
rect 3850 34644 4260 34647
rect 5031 34638 5034 34696
rect 5060 34638 5063 34696
rect 5031 34635 5063 34638
rect 5090 34618 5170 34925
rect 14790 34967 14870 35325
rect 16233 35242 16283 35245
rect 16233 35198 16236 35242
rect 16280 35198 16283 35242
rect 16233 35195 16283 35198
rect 14913 35187 14971 35190
rect 14913 35135 14916 35187
rect 14968 35135 14971 35187
rect 14913 35132 14971 35135
rect 16233 35178 16283 35181
rect 16233 35134 16236 35178
rect 16280 35134 16283 35178
rect 16233 35131 16283 35134
rect 14897 35096 14929 35099
rect 14897 35038 14900 35096
rect 14926 35038 14929 35096
rect 15700 35047 15703 35073
rect 16107 35047 16110 35073
rect 15700 35042 16110 35047
rect 14897 35035 14929 35038
rect 16718 35007 16768 39198
rect 14790 34925 16287 34967
rect 16718 34949 16721 35007
rect 16765 34949 16768 35007
rect 16718 34946 16768 34949
rect 16782 39192 16832 39195
rect 16782 39134 16785 39192
rect 16829 39134 16832 39192
rect 14790 34618 14870 34925
rect 16782 34917 16832 39134
rect 16782 34859 16785 34917
rect 16829 34859 16832 34917
rect 16782 34856 16832 34859
rect 16846 38856 16896 38859
rect 16846 38798 16849 38856
rect 16893 38798 16896 38856
rect 16233 34842 16283 34845
rect 16233 34798 16236 34842
rect 16280 34798 16283 34842
rect 16233 34795 16283 34798
rect 14913 34787 14971 34790
rect 14913 34735 14916 34787
rect 14968 34735 14971 34787
rect 14913 34732 14971 34735
rect 16233 34778 16283 34781
rect 16233 34734 16236 34778
rect 16280 34734 16283 34778
rect 16233 34731 16283 34734
rect 14897 34696 14929 34699
rect 14897 34638 14900 34696
rect 14926 34638 14929 34696
rect 15700 34647 15703 34673
rect 16107 34647 16110 34673
rect 15700 34642 16110 34647
rect 14897 34635 14929 34638
rect 5090 34567 5141 34618
rect 3673 34560 5141 34567
rect 5167 34560 5170 34618
rect 14790 34560 14793 34618
rect 14819 34567 14870 34618
rect 14819 34560 16287 34567
rect 3673 34525 5170 34560
rect 3677 34442 3727 34445
rect 3677 34398 3680 34442
rect 3724 34398 3727 34442
rect 3677 34395 3727 34398
rect 4989 34387 5047 34390
rect 3677 34378 3727 34381
rect 3677 34334 3680 34378
rect 3724 34334 3727 34378
rect 3677 34331 3727 34334
rect 4989 34335 4992 34387
rect 5044 34335 5047 34387
rect 4989 34332 5047 34335
rect 5031 34296 5063 34299
rect 3850 34247 3853 34273
rect 4257 34247 4260 34273
rect 3850 34244 4260 34247
rect 5031 34238 5034 34296
rect 5060 34238 5063 34296
rect 5031 34235 5063 34238
rect 5090 34167 5170 34525
rect 14790 34525 16287 34560
rect 3673 34125 5170 34167
rect 3677 34042 3727 34045
rect 3677 33998 3680 34042
rect 3724 33998 3727 34042
rect 3677 33995 3727 33998
rect 4989 33987 5047 33990
rect 3677 33978 3727 33981
rect 3677 33934 3680 33978
rect 3724 33934 3727 33978
rect 3677 33931 3727 33934
rect 4989 33935 4992 33987
rect 5044 33935 5047 33987
rect 4989 33932 5047 33935
rect 5031 33896 5063 33899
rect 3850 33847 3853 33873
rect 4257 33847 4260 33873
rect 3850 33844 4260 33847
rect 5031 33838 5034 33896
rect 5060 33838 5063 33896
rect 5031 33835 5063 33838
rect 5090 33818 5170 34125
rect 14790 34167 14870 34525
rect 16233 34442 16283 34445
rect 16233 34398 16236 34442
rect 16280 34398 16283 34442
rect 16233 34395 16283 34398
rect 14913 34387 14971 34390
rect 14913 34335 14916 34387
rect 14968 34335 14971 34387
rect 14913 34332 14971 34335
rect 16233 34378 16283 34381
rect 16233 34334 16236 34378
rect 16280 34334 16283 34378
rect 16233 34331 16283 34334
rect 14897 34296 14929 34299
rect 14897 34238 14900 34296
rect 14926 34238 14929 34296
rect 15700 34247 15703 34273
rect 16107 34247 16110 34273
rect 15700 34242 16110 34247
rect 14897 34235 14929 34238
rect 14790 34125 16287 34167
rect 14790 33818 14870 34125
rect 16233 34042 16283 34045
rect 16233 33998 16236 34042
rect 16280 33998 16283 34042
rect 16233 33995 16283 33998
rect 14913 33987 14971 33990
rect 14913 33935 14916 33987
rect 14968 33935 14971 33987
rect 14913 33932 14971 33935
rect 16233 33978 16283 33981
rect 16233 33934 16236 33978
rect 16280 33934 16283 33978
rect 16233 33931 16283 33934
rect 14897 33896 14929 33899
rect 14897 33838 14900 33896
rect 14926 33838 14929 33896
rect 15700 33847 15703 33873
rect 16107 33847 16110 33873
rect 15700 33842 16110 33847
rect 14897 33835 14929 33838
rect 5090 33767 5141 33818
rect 3673 33760 5141 33767
rect 5167 33760 5170 33818
rect 14790 33760 14793 33818
rect 14819 33767 14870 33818
rect 14819 33760 16287 33767
rect 3673 33725 5170 33760
rect 3677 33642 3727 33645
rect 3677 33598 3680 33642
rect 3724 33598 3727 33642
rect 3677 33595 3727 33598
rect 4989 33587 5047 33590
rect 3677 33578 3727 33581
rect 3677 33534 3680 33578
rect 3724 33534 3727 33578
rect 3677 33531 3727 33534
rect 4989 33535 4992 33587
rect 5044 33535 5047 33587
rect 4989 33532 5047 33535
rect 3064 33449 3067 33507
rect 3111 33449 3114 33507
rect 5031 33496 5063 33499
rect 3064 33446 3114 33449
rect 3850 33447 3853 33473
rect 4257 33447 4260 33473
rect 3850 33444 4260 33447
rect 5031 33438 5034 33496
rect 5060 33438 5063 33496
rect 5031 33435 5063 33438
rect 3000 33359 3003 33417
rect 3047 33359 3050 33417
rect 5090 33367 5170 33725
rect 14790 33725 16287 33760
rect 3000 33356 3050 33359
rect 3673 33325 5170 33367
rect 3677 33242 3727 33245
rect 3677 33198 3680 33242
rect 3724 33198 3727 33242
rect 3677 33195 3727 33198
rect 4989 33187 5047 33190
rect 3677 33178 3727 33181
rect 3677 33134 3680 33178
rect 3724 33134 3727 33178
rect 3677 33131 3727 33134
rect 4989 33135 4992 33187
rect 5044 33135 5047 33187
rect 4989 33132 5047 33135
rect 5031 33096 5063 33099
rect 3850 33047 3853 33073
rect 4257 33047 4260 33073
rect 3850 33044 4260 33047
rect 5031 33038 5034 33096
rect 5060 33038 5063 33096
rect 5031 33035 5063 33038
rect 5090 33018 5170 33325
rect 14790 33367 14870 33725
rect 16233 33642 16283 33645
rect 16233 33598 16236 33642
rect 16280 33598 16283 33642
rect 16233 33595 16283 33598
rect 14913 33587 14971 33590
rect 14913 33535 14916 33587
rect 14968 33535 14971 33587
rect 14913 33532 14971 33535
rect 16233 33578 16283 33581
rect 16233 33534 16236 33578
rect 16280 33534 16283 33578
rect 16233 33531 16283 33534
rect 16846 33507 16896 38798
rect 14897 33496 14929 33499
rect 14897 33438 14900 33496
rect 14926 33438 14929 33496
rect 15700 33447 15703 33473
rect 16107 33447 16110 33473
rect 15700 33442 16110 33447
rect 16846 33449 16849 33507
rect 16893 33449 16896 33507
rect 16846 33446 16896 33449
rect 16910 38792 16960 38795
rect 16910 38734 16913 38792
rect 16957 38734 16960 38792
rect 14897 33435 14929 33438
rect 16910 33417 16960 38734
rect 14790 33325 16287 33367
rect 16910 33359 16913 33417
rect 16957 33359 16960 33417
rect 16910 33356 16960 33359
rect 16974 38456 17024 38459
rect 16974 38398 16977 38456
rect 17021 38398 17024 38456
rect 14790 33018 14870 33325
rect 16233 33242 16283 33245
rect 16233 33198 16236 33242
rect 16280 33198 16283 33242
rect 16233 33195 16283 33198
rect 14913 33187 14971 33190
rect 14913 33135 14916 33187
rect 14968 33135 14971 33187
rect 14913 33132 14971 33135
rect 16233 33178 16283 33181
rect 16233 33134 16236 33178
rect 16280 33134 16283 33178
rect 16233 33131 16283 33134
rect 14897 33096 14929 33099
rect 14897 33038 14900 33096
rect 14926 33038 14929 33096
rect 15700 33047 15703 33073
rect 16107 33047 16110 33073
rect 15700 33042 16110 33047
rect 14897 33035 14929 33038
rect 5090 32967 5141 33018
rect 3673 32960 5141 32967
rect 5167 32960 5170 33018
rect 14790 32960 14793 33018
rect 14819 32967 14870 33018
rect 14819 32960 16287 32967
rect 3673 32925 5170 32960
rect 3677 32842 3727 32845
rect 3677 32798 3680 32842
rect 3724 32798 3727 32842
rect 3677 32795 3727 32798
rect 4989 32787 5047 32790
rect 3677 32778 3727 32781
rect 3677 32734 3680 32778
rect 3724 32734 3727 32778
rect 3677 32731 3727 32734
rect 4989 32735 4992 32787
rect 5044 32735 5047 32787
rect 4989 32732 5047 32735
rect 5031 32696 5063 32699
rect 3850 32647 3853 32673
rect 4257 32647 4260 32673
rect 3850 32644 4260 32647
rect 5031 32638 5034 32696
rect 5060 32638 5063 32696
rect 5031 32635 5063 32638
rect 5090 32567 5170 32925
rect 14790 32925 16287 32960
rect 3673 32525 5170 32567
rect 3677 32442 3727 32445
rect 3677 32398 3680 32442
rect 3724 32398 3727 32442
rect 3677 32395 3727 32398
rect 4989 32387 5047 32390
rect 3677 32378 3727 32381
rect 3677 32334 3680 32378
rect 3724 32334 3727 32378
rect 3677 32331 3727 32334
rect 4989 32335 4992 32387
rect 5044 32335 5047 32387
rect 4989 32332 5047 32335
rect 5031 32296 5063 32299
rect 3850 32247 3853 32273
rect 4257 32247 4260 32273
rect 3850 32244 4260 32247
rect 5031 32238 5034 32296
rect 5060 32238 5063 32296
rect 5031 32235 5063 32238
rect 5090 32218 5170 32525
rect 14790 32567 14870 32925
rect 16233 32842 16283 32845
rect 16233 32798 16236 32842
rect 16280 32798 16283 32842
rect 16233 32795 16283 32798
rect 14913 32787 14971 32790
rect 14913 32735 14916 32787
rect 14968 32735 14971 32787
rect 14913 32732 14971 32735
rect 16233 32778 16283 32781
rect 16233 32734 16236 32778
rect 16280 32734 16283 32778
rect 16233 32731 16283 32734
rect 14897 32696 14929 32699
rect 14897 32638 14900 32696
rect 14926 32638 14929 32696
rect 15700 32647 15703 32673
rect 16107 32647 16110 32673
rect 15700 32642 16110 32647
rect 14897 32635 14929 32638
rect 14790 32525 16287 32567
rect 14790 32218 14870 32525
rect 16233 32442 16283 32445
rect 16233 32398 16236 32442
rect 16280 32398 16283 32442
rect 16233 32395 16283 32398
rect 14913 32387 14971 32390
rect 14913 32335 14916 32387
rect 14968 32335 14971 32387
rect 14913 32332 14971 32335
rect 16233 32378 16283 32381
rect 16233 32334 16236 32378
rect 16280 32334 16283 32378
rect 16233 32331 16283 32334
rect 14897 32296 14929 32299
rect 14897 32238 14900 32296
rect 14926 32238 14929 32296
rect 15700 32247 15703 32273
rect 16107 32247 16110 32273
rect 15700 32242 16110 32247
rect 14897 32235 14929 32238
rect 5090 32167 5141 32218
rect 3673 32160 5141 32167
rect 5167 32160 5170 32218
rect 14790 32160 14793 32218
rect 14819 32167 14870 32218
rect 14819 32160 16287 32167
rect 3673 32125 5170 32160
rect 2936 31949 2939 32007
rect 2983 31949 2986 32007
rect 3677 32042 3727 32045
rect 3677 31998 3680 32042
rect 3724 31998 3727 32042
rect 3677 31995 3727 31998
rect 4989 31987 5047 31990
rect 2936 31946 2986 31949
rect 3677 31978 3727 31981
rect 3677 31934 3680 31978
rect 3724 31934 3727 31978
rect 3677 31931 3727 31934
rect 4989 31935 4992 31987
rect 5044 31935 5047 31987
rect 4989 31932 5047 31935
rect 2872 31859 2875 31917
rect 2919 31859 2922 31917
rect 5031 31896 5063 31899
rect 2872 31856 2922 31859
rect 3850 31847 3853 31873
rect 4257 31847 4260 31873
rect 3850 31844 4260 31847
rect 5031 31838 5034 31896
rect 5060 31838 5063 31896
rect 5031 31835 5063 31838
rect 5090 31767 5170 32125
rect 14790 32125 16287 32160
rect 3673 31725 5170 31767
rect 3677 31642 3727 31645
rect 3677 31598 3680 31642
rect 3724 31598 3727 31642
rect 3677 31595 3727 31598
rect 4989 31587 5047 31590
rect 3677 31578 3727 31581
rect 3677 31534 3680 31578
rect 3724 31534 3727 31578
rect 3677 31531 3727 31534
rect 4989 31535 4992 31587
rect 5044 31535 5047 31587
rect 4989 31532 5047 31535
rect 5031 31496 5063 31499
rect 3850 31447 3853 31473
rect 4257 31447 4260 31473
rect 3850 31444 4260 31447
rect 5031 31438 5034 31496
rect 5060 31438 5063 31496
rect 5031 31435 5063 31438
rect 5090 31418 5170 31725
rect 14790 31767 14870 32125
rect 16233 32042 16283 32045
rect 16233 31998 16236 32042
rect 16280 31998 16283 32042
rect 16233 31995 16283 31998
rect 16974 32007 17024 38398
rect 14913 31987 14971 31990
rect 14913 31935 14916 31987
rect 14968 31935 14971 31987
rect 14913 31932 14971 31935
rect 16233 31978 16283 31981
rect 16233 31934 16236 31978
rect 16280 31934 16283 31978
rect 16974 31949 16977 32007
rect 17021 31949 17024 32007
rect 16974 31946 17024 31949
rect 17038 38392 17088 38395
rect 17038 38334 17041 38392
rect 17085 38334 17088 38392
rect 16233 31931 16283 31934
rect 17038 31917 17088 38334
rect 14897 31896 14929 31899
rect 14897 31838 14900 31896
rect 14926 31838 14929 31896
rect 15700 31847 15703 31873
rect 16107 31847 16110 31873
rect 17038 31859 17041 31917
rect 17085 31859 17088 31917
rect 17038 31856 17088 31859
rect 17102 38155 17152 38158
rect 17102 38097 17105 38155
rect 17149 38097 17152 38155
rect 15700 31842 16110 31847
rect 14897 31835 14929 31838
rect 14790 31725 16287 31767
rect 14790 31418 14870 31725
rect 16233 31642 16283 31645
rect 16233 31598 16236 31642
rect 16280 31598 16283 31642
rect 16233 31595 16283 31598
rect 14913 31587 14971 31590
rect 14913 31535 14916 31587
rect 14968 31535 14971 31587
rect 14913 31532 14971 31535
rect 16233 31578 16283 31581
rect 16233 31534 16236 31578
rect 16280 31534 16283 31578
rect 16233 31531 16283 31534
rect 14897 31496 14929 31499
rect 14897 31438 14900 31496
rect 14926 31438 14929 31496
rect 15700 31447 15703 31473
rect 16107 31447 16110 31473
rect 15700 31442 16110 31447
rect 14897 31435 14929 31438
rect 5090 31367 5141 31418
rect 3673 31360 5141 31367
rect 5167 31360 5170 31418
rect 14790 31360 14793 31418
rect 14819 31367 14870 31418
rect 14819 31360 16287 31367
rect 3673 31325 5170 31360
rect 3677 31242 3727 31245
rect 3677 31198 3680 31242
rect 3724 31198 3727 31242
rect 3677 31195 3727 31198
rect 4989 31187 5047 31190
rect 3677 31178 3727 31181
rect 3677 31134 3680 31178
rect 3724 31134 3727 31178
rect 3677 31131 3727 31134
rect 4989 31135 4992 31187
rect 5044 31135 5047 31187
rect 4989 31132 5047 31135
rect 5031 31096 5063 31099
rect 3850 31047 3853 31073
rect 4257 31047 4260 31073
rect 3850 31044 4260 31047
rect 5031 31038 5034 31096
rect 5060 31038 5063 31096
rect 5031 31035 5063 31038
rect 5090 30967 5170 31325
rect 14790 31325 16287 31360
rect 3673 30925 5170 30967
rect 3677 30842 3727 30845
rect 3677 30798 3680 30842
rect 3724 30798 3727 30842
rect 3677 30795 3727 30798
rect 4989 30787 5047 30790
rect 3677 30778 3727 30781
rect 3677 30734 3680 30778
rect 3724 30734 3727 30778
rect 3677 30731 3727 30734
rect 4989 30735 4992 30787
rect 5044 30735 5047 30787
rect 4989 30732 5047 30735
rect 5031 30696 5063 30699
rect 3850 30647 3853 30673
rect 4257 30647 4260 30673
rect 3850 30644 4260 30647
rect 5031 30638 5034 30696
rect 5060 30638 5063 30696
rect 5031 30635 5063 30638
rect 5090 30618 5170 30925
rect 14790 30967 14870 31325
rect 16233 31242 16283 31245
rect 16233 31198 16236 31242
rect 16280 31198 16283 31242
rect 16233 31195 16283 31198
rect 14913 31187 14971 31190
rect 14913 31135 14916 31187
rect 14968 31135 14971 31187
rect 14913 31132 14971 31135
rect 16233 31178 16283 31181
rect 16233 31134 16236 31178
rect 16280 31134 16283 31178
rect 16233 31131 16283 31134
rect 14897 31096 14929 31099
rect 14897 31038 14900 31096
rect 14926 31038 14929 31096
rect 15700 31047 15703 31073
rect 16107 31047 16110 31073
rect 15700 31042 16110 31047
rect 14897 31035 14929 31038
rect 14790 30925 16287 30967
rect 14790 30618 14870 30925
rect 16233 30842 16283 30845
rect 16233 30798 16236 30842
rect 16280 30798 16283 30842
rect 16233 30795 16283 30798
rect 14913 30787 14971 30790
rect 14913 30735 14916 30787
rect 14968 30735 14971 30787
rect 14913 30732 14971 30735
rect 16233 30778 16283 30781
rect 16233 30734 16236 30778
rect 16280 30734 16283 30778
rect 16233 30731 16283 30734
rect 14897 30696 14929 30699
rect 14897 30638 14900 30696
rect 14926 30638 14929 30696
rect 15700 30647 15703 30673
rect 16107 30647 16110 30673
rect 15700 30642 16110 30647
rect 14897 30635 14929 30638
rect 5090 30567 5141 30618
rect 3673 30560 5141 30567
rect 5167 30560 5170 30618
rect 14790 30560 14793 30618
rect 14819 30567 14870 30618
rect 14819 30560 16287 30567
rect 3673 30525 5170 30560
rect 2808 30449 2811 30507
rect 2855 30449 2858 30507
rect 2808 30446 2858 30449
rect 2744 30359 2747 30417
rect 2791 30359 2794 30417
rect 3677 30442 3727 30445
rect 3677 30398 3680 30442
rect 3724 30398 3727 30442
rect 3677 30395 3727 30398
rect 4989 30387 5047 30390
rect 2744 30356 2794 30359
rect 3677 30378 3727 30381
rect 3677 30334 3680 30378
rect 3724 30334 3727 30378
rect 3677 30331 3727 30334
rect 4989 30335 4992 30387
rect 5044 30335 5047 30387
rect 4989 30332 5047 30335
rect 5031 30296 5063 30299
rect 3850 30247 3853 30273
rect 4257 30247 4260 30273
rect 3850 30244 4260 30247
rect 5031 30238 5034 30296
rect 5060 30238 5063 30296
rect 5031 30235 5063 30238
rect 5090 30167 5170 30525
rect 14790 30525 16287 30560
rect 3673 30125 5170 30167
rect 3677 30042 3727 30045
rect 3677 29998 3680 30042
rect 3724 29998 3727 30042
rect 3677 29995 3727 29998
rect 4989 29987 5047 29990
rect 3677 29978 3727 29981
rect 3677 29934 3680 29978
rect 3724 29934 3727 29978
rect 3677 29931 3727 29934
rect 4989 29935 4992 29987
rect 5044 29935 5047 29987
rect 4989 29932 5047 29935
rect 5031 29896 5063 29899
rect 3850 29847 3853 29873
rect 4257 29847 4260 29873
rect 3850 29844 4260 29847
rect 5031 29838 5034 29896
rect 5060 29838 5063 29896
rect 5031 29835 5063 29838
rect 5090 29818 5170 30125
rect 14790 30167 14870 30525
rect 17102 30507 17152 38097
rect 17102 30449 17105 30507
rect 17149 30449 17152 30507
rect 17102 30446 17152 30449
rect 17166 38091 17216 38094
rect 17166 38033 17169 38091
rect 17213 38033 17216 38091
rect 16233 30442 16283 30445
rect 16233 30398 16236 30442
rect 16280 30398 16283 30442
rect 16233 30395 16283 30398
rect 17166 30417 17216 38033
rect 14913 30387 14971 30390
rect 14913 30335 14916 30387
rect 14968 30335 14971 30387
rect 14913 30332 14971 30335
rect 16233 30378 16283 30381
rect 16233 30334 16236 30378
rect 16280 30334 16283 30378
rect 17166 30359 17169 30417
rect 17213 30359 17216 30417
rect 17166 30356 17216 30359
rect 17230 37656 17280 37659
rect 17230 37598 17233 37656
rect 17277 37598 17280 37656
rect 16233 30331 16283 30334
rect 14897 30296 14929 30299
rect 14897 30238 14900 30296
rect 14926 30238 14929 30296
rect 15700 30247 15703 30273
rect 16107 30247 16110 30273
rect 15700 30242 16110 30247
rect 14897 30235 14929 30238
rect 14790 30125 16287 30167
rect 14790 29818 14870 30125
rect 16233 30042 16283 30045
rect 16233 29998 16236 30042
rect 16280 29998 16283 30042
rect 16233 29995 16283 29998
rect 14913 29987 14971 29990
rect 14913 29935 14916 29987
rect 14968 29935 14971 29987
rect 14913 29932 14971 29935
rect 16233 29978 16283 29981
rect 16233 29934 16236 29978
rect 16280 29934 16283 29978
rect 16233 29931 16283 29934
rect 14897 29896 14929 29899
rect 14897 29838 14900 29896
rect 14926 29838 14929 29896
rect 15700 29847 15703 29873
rect 16107 29847 16110 29873
rect 15700 29842 16110 29847
rect 14897 29835 14929 29838
rect 5090 29767 5141 29818
rect 3673 29760 5141 29767
rect 5167 29760 5170 29818
rect 14790 29760 14793 29818
rect 14819 29767 14870 29818
rect 14819 29760 16287 29767
rect 3673 29725 5170 29760
rect 3677 29642 3727 29645
rect 3677 29598 3680 29642
rect 3724 29598 3727 29642
rect 3677 29595 3727 29598
rect 4989 29587 5047 29590
rect 3677 29578 3727 29581
rect 3677 29534 3680 29578
rect 3724 29534 3727 29578
rect 3677 29531 3727 29534
rect 4989 29535 4992 29587
rect 5044 29535 5047 29587
rect 4989 29532 5047 29535
rect 5031 29496 5063 29499
rect 3850 29447 3853 29473
rect 4257 29447 4260 29473
rect 3850 29444 4260 29447
rect 5031 29438 5034 29496
rect 5060 29438 5063 29496
rect 5031 29435 5063 29438
rect 5090 29367 5170 29725
rect 14790 29725 16287 29760
rect 3673 29325 5170 29367
rect 14790 29367 14870 29725
rect 16233 29642 16283 29645
rect 16233 29598 16236 29642
rect 16280 29598 16283 29642
rect 16233 29595 16283 29598
rect 14913 29587 14971 29590
rect 14913 29535 14916 29587
rect 14968 29535 14971 29587
rect 14913 29532 14971 29535
rect 16233 29578 16283 29581
rect 16233 29534 16236 29578
rect 16280 29534 16283 29578
rect 16233 29531 16283 29534
rect 14897 29496 14929 29499
rect 14897 29438 14900 29496
rect 14926 29438 14929 29496
rect 15700 29447 15703 29473
rect 16107 29447 16110 29473
rect 15700 29442 16110 29447
rect 14897 29435 14929 29438
rect 3677 29242 3727 29245
rect 3677 29198 3680 29242
rect 3724 29198 3727 29242
rect 3677 29195 3727 29198
rect 4989 29187 5047 29190
rect 3677 29178 3727 29181
rect 3677 29134 3680 29178
rect 3724 29134 3727 29178
rect 3677 29131 3727 29134
rect 4989 29135 4992 29187
rect 5044 29135 5047 29187
rect 4989 29132 5047 29135
rect 5031 29096 5063 29099
rect 3850 29047 3853 29073
rect 4257 29047 4260 29073
rect 3850 29044 4260 29047
rect 5031 29038 5034 29096
rect 5060 29038 5063 29096
rect 5031 29035 5063 29038
rect 2680 28949 2683 29007
rect 2727 28949 2730 29007
rect 2680 28946 2730 28949
rect 5090 29000 5170 29325
rect 5210 29096 5290 29352
rect 5210 29038 5213 29096
rect 5239 29038 5290 29096
rect 5210 29035 5290 29038
rect 14670 29096 14750 29353
rect 14670 29038 14721 29096
rect 14747 29038 14750 29096
rect 14670 29035 14750 29038
rect 14790 29325 16287 29367
rect 14790 29000 14870 29325
rect 16233 29242 16283 29245
rect 16233 29198 16236 29242
rect 16280 29198 16283 29242
rect 16233 29195 16283 29198
rect 14913 29187 14971 29190
rect 14913 29135 14916 29187
rect 14968 29135 14971 29187
rect 14913 29132 14971 29135
rect 16233 29178 16283 29181
rect 16233 29134 16236 29178
rect 16280 29134 16283 29178
rect 16233 29131 16283 29134
rect 14897 29096 14929 29099
rect 14897 29038 14900 29096
rect 14926 29038 14929 29096
rect 15700 29047 15703 29073
rect 16107 29047 16110 29073
rect 15700 29042 16110 29047
rect 14897 29035 14929 29038
rect 5090 28997 5820 29000
rect 2616 28859 2619 28917
rect 2663 28859 2666 28917
rect 5090 28908 5175 28997
rect 5815 28908 5820 28997
rect 5090 28903 5820 28908
rect 14140 28997 14870 29000
rect 14140 28908 14145 28997
rect 14785 28908 14870 28997
rect 17230 29007 17280 37598
rect 17230 28949 17233 29007
rect 17277 28949 17280 29007
rect 17230 28946 17280 28949
rect 17294 37592 17344 37595
rect 17294 37534 17297 37592
rect 17341 37534 17344 37592
rect 14140 28903 14870 28908
rect 17294 28917 17344 37534
rect 2616 28856 2666 28859
rect 17294 28859 17297 28917
rect 17341 28859 17344 28917
rect 17294 28856 17344 28859
rect 17358 37256 17408 37259
rect 17358 37198 17361 37256
rect 17405 37198 17408 37256
rect 2552 27449 2555 27507
rect 2599 27449 2602 27507
rect 2552 27446 2602 27449
rect 17358 27507 17408 37198
rect 17358 27449 17361 27507
rect 17405 27449 17408 27507
rect 17358 27446 17408 27449
rect 17422 37192 17472 37195
rect 17422 37134 17425 37192
rect 17469 37134 17472 37192
rect 2488 27359 2491 27417
rect 2535 27359 2538 27417
rect 2488 27356 2538 27359
rect 17422 27417 17472 37134
rect 17422 27359 17425 27417
rect 17469 27359 17472 27417
rect 17422 27356 17472 27359
rect 17486 36856 17536 36859
rect 17486 36798 17489 36856
rect 17533 36798 17536 36856
rect 2424 25949 2427 26007
rect 2471 25949 2474 26007
rect 2424 25946 2474 25949
rect 17486 26007 17536 36798
rect 17486 25949 17489 26007
rect 17533 25949 17536 26007
rect 17486 25946 17536 25949
rect 17550 36792 17600 36795
rect 17550 36734 17553 36792
rect 17597 36734 17600 36792
rect 2360 25859 2363 25917
rect 2407 25859 2410 25917
rect 2360 25856 2410 25859
rect 17550 25917 17600 36734
rect 17550 25859 17553 25917
rect 17597 25859 17600 25917
rect 17550 25856 17600 25859
rect 17614 36655 17664 36658
rect 17614 36597 17617 36655
rect 17661 36597 17664 36655
rect 2296 24449 2299 24507
rect 2343 24449 2346 24507
rect 2296 24446 2346 24449
rect 17614 24507 17664 36597
rect 17614 24449 17617 24507
rect 17661 24449 17664 24507
rect 17614 24446 17664 24449
rect 17678 36591 17728 36594
rect 17678 36533 17681 36591
rect 17725 36533 17728 36591
rect 2232 24359 2235 24417
rect 2279 24359 2282 24417
rect 2232 24356 2282 24359
rect 17678 24417 17728 36533
rect 17678 24359 17681 24417
rect 17725 24359 17728 24417
rect 17678 24356 17728 24359
rect 17742 36056 17792 36059
rect 17742 35998 17745 36056
rect 17789 35998 17792 36056
rect 2168 22949 2171 23007
rect 2215 22949 2218 23007
rect 2168 22946 2218 22949
rect 17742 23007 17792 35998
rect 17742 22949 17745 23007
rect 17789 22949 17792 23007
rect 17742 22946 17792 22949
rect 17806 35992 17856 35995
rect 17806 35934 17809 35992
rect 17853 35934 17856 35992
rect 2104 22859 2107 22917
rect 2151 22859 2154 22917
rect 2104 22856 2154 22859
rect 17806 22917 17856 35934
rect 17806 22859 17809 22917
rect 17853 22859 17856 22917
rect 17806 22856 17856 22859
rect 17870 35656 17920 35659
rect 17870 35598 17873 35656
rect 17917 35598 17920 35656
rect 2040 21449 2043 21507
rect 2087 21449 2090 21507
rect 2040 21446 2090 21449
rect 17870 21507 17920 35598
rect 17870 21449 17873 21507
rect 17917 21449 17920 21507
rect 17870 21446 17920 21449
rect 17934 35592 17984 35595
rect 17934 35534 17937 35592
rect 17981 35534 17984 35592
rect 1976 21359 1979 21417
rect 2023 21359 2026 21417
rect 1976 21356 2026 21359
rect 17934 21417 17984 35534
rect 17934 21359 17937 21417
rect 17981 21359 17984 21417
rect 17934 21356 17984 21359
rect 17998 35256 18048 35259
rect 17998 35198 18001 35256
rect 18045 35198 18048 35256
rect 3300 21295 5820 21300
rect 3300 21105 5175 21295
rect 5815 21105 5820 21295
rect 3300 21100 5820 21105
rect 14140 21295 16541 21300
rect 14140 21105 14145 21295
rect 14785 21105 16541 21295
rect 14140 21100 16541 21105
rect 3300 21087 4441 21100
rect 3300 21070 3312 21087
rect 4428 21070 4441 21087
rect 3300 21069 4441 21070
rect 15400 21089 16541 21100
rect 15400 21072 15412 21089
rect 16528 21072 16541 21089
rect 15400 21069 16541 21072
rect 1912 19949 1915 20007
rect 1959 19949 1962 20007
rect 1912 19946 1962 19949
rect 17998 20007 18048 35198
rect 17998 19949 18001 20007
rect 18045 19949 18048 20007
rect 17998 19946 18048 19949
rect 18062 35192 18112 35195
rect 18062 35134 18065 35192
rect 18109 35134 18112 35192
rect 1848 19859 1851 19917
rect 1895 19859 1898 19917
rect 1848 19856 1898 19859
rect 18062 19917 18112 35134
rect 18062 19859 18065 19917
rect 18109 19859 18112 19917
rect 18062 19856 18112 19859
rect 18126 34853 18176 34856
rect 18126 34795 18129 34853
rect 18173 34795 18176 34853
rect 10965 19460 11095 19465
rect 10965 19340 10970 19460
rect 11090 19340 11095 19460
rect 10965 19335 11095 19340
rect 10590 19277 10649 19280
rect 10590 19066 10593 19277
rect 10646 19066 10649 19277
rect 11114 19273 11174 19276
rect 10590 19063 10649 19066
rect 10999 19270 11040 19273
rect 10999 19060 11002 19270
rect 11037 19060 11040 19270
rect 11114 19063 11117 19273
rect 11171 19063 11174 19273
rect 11114 19060 11174 19063
rect 10999 19057 11040 19060
rect 1784 18449 1787 18507
rect 1831 18449 1834 18507
rect 1784 18446 1834 18449
rect 18126 18507 18176 34795
rect 18126 18449 18129 18507
rect 18173 18449 18176 18507
rect 18126 18446 18176 18449
rect 18190 34789 18240 34792
rect 18190 34731 18193 34789
rect 18237 34731 18240 34789
rect 1720 18359 1723 18417
rect 1767 18359 1770 18417
rect 1720 18356 1770 18359
rect 18190 18417 18240 34731
rect 18190 18359 18193 18417
rect 18237 18359 18240 18417
rect 18190 18356 18240 18359
rect 18254 34456 18304 34459
rect 18254 34398 18257 34456
rect 18301 34398 18304 34456
rect 1656 16949 1659 17007
rect 1703 16949 1706 17007
rect 1656 16946 1706 16949
rect 18254 17007 18304 34398
rect 18254 16949 18257 17007
rect 18301 16949 18304 17007
rect 18254 16946 18304 16949
rect 18318 34392 18368 34395
rect 18318 34334 18321 34392
rect 18365 34334 18368 34392
rect 1592 16859 1595 16917
rect 1639 16859 1642 16917
rect 1592 16856 1642 16859
rect 18318 16917 18368 34334
rect 18318 16859 18321 16917
rect 18365 16859 18368 16917
rect 18318 16856 18368 16859
rect 18382 34056 18432 34059
rect 18382 33998 18385 34056
rect 18429 33998 18432 34056
rect 1528 15449 1531 15507
rect 1575 15449 1578 15507
rect 1528 15446 1578 15449
rect 18382 15507 18432 33998
rect 18382 15449 18385 15507
rect 18429 15449 18432 15507
rect 18382 15446 18432 15449
rect 18446 33992 18496 33995
rect 18446 33934 18449 33992
rect 18493 33934 18496 33992
rect 1464 15359 1467 15417
rect 1511 15359 1514 15417
rect 1464 15356 1514 15359
rect 18446 15417 18496 33934
rect 18446 15359 18449 15417
rect 18493 15359 18496 15417
rect 18446 15356 18496 15359
rect 18510 33656 18560 33659
rect 18510 33598 18513 33656
rect 18557 33598 18560 33656
rect 1400 13949 1403 14007
rect 1447 13949 1450 14007
rect 1400 13946 1450 13949
rect 18510 14007 18560 33598
rect 18510 13949 18513 14007
rect 18557 13949 18560 14007
rect 18510 13946 18560 13949
rect 18574 33592 18624 33595
rect 18574 33534 18577 33592
rect 18621 33534 18624 33592
rect 1336 13859 1339 13917
rect 1383 13859 1386 13917
rect 1336 13856 1386 13859
rect 18574 13917 18624 33534
rect 18574 13859 18577 13917
rect 18621 13859 18624 13917
rect 18574 13856 18624 13859
rect 18638 33256 18688 33259
rect 18638 33198 18641 33256
rect 18685 33198 18688 33256
rect 1272 12449 1275 12507
rect 1319 12449 1322 12507
rect 1272 12446 1322 12449
rect 18638 12507 18688 33198
rect 18638 12449 18641 12507
rect 18685 12449 18688 12507
rect 18638 12446 18688 12449
rect 18702 33192 18752 33195
rect 18702 33134 18705 33192
rect 18749 33134 18752 33192
rect 1208 12359 1211 12417
rect 1255 12359 1258 12417
rect 1208 12356 1258 12359
rect 18702 12417 18752 33134
rect 18702 12359 18705 12417
rect 18749 12359 18752 12417
rect 18702 12356 18752 12359
rect 18766 32856 18816 32859
rect 18766 32798 18769 32856
rect 18813 32798 18816 32856
rect 1144 10949 1147 11007
rect 1191 10949 1194 11007
rect 1144 10946 1194 10949
rect 18766 11007 18816 32798
rect 18766 10949 18769 11007
rect 18813 10949 18816 11007
rect 18766 10946 18816 10949
rect 18830 32792 18880 32795
rect 18830 32734 18833 32792
rect 18877 32734 18880 32792
rect 1080 10859 1083 10917
rect 1127 10859 1130 10917
rect 1080 10856 1130 10859
rect 18830 10917 18880 32734
rect 18830 10859 18833 10917
rect 18877 10859 18880 10917
rect 18830 10856 18880 10859
rect 18894 32456 18944 32459
rect 18894 32398 18897 32456
rect 18941 32398 18944 32456
rect 1016 9449 1019 9507
rect 1063 9449 1066 9507
rect 1016 9446 1066 9449
rect 18894 9507 18944 32398
rect 18894 9449 18897 9507
rect 18941 9449 18944 9507
rect 18894 9446 18944 9449
rect 18958 32392 19008 32395
rect 18958 32334 18961 32392
rect 19005 32334 19008 32392
rect 952 9359 955 9417
rect 999 9359 1002 9417
rect 952 9356 1002 9359
rect 18958 9417 19008 32334
rect 18958 9359 18961 9417
rect 19005 9359 19008 9417
rect 18958 9356 19008 9359
rect 19022 32149 19072 32152
rect 19022 32091 19025 32149
rect 19069 32091 19072 32149
rect 888 7949 891 8007
rect 935 7949 938 8007
rect 888 7946 938 7949
rect 19022 8007 19072 32091
rect 19022 7949 19025 8007
rect 19069 7949 19072 8007
rect 19022 7946 19072 7949
rect 19086 32085 19136 32088
rect 19086 32027 19089 32085
rect 19133 32027 19136 32085
rect 824 7859 827 7917
rect 871 7859 874 7917
rect 824 7856 874 7859
rect 19086 7917 19136 32027
rect 19086 7859 19089 7917
rect 19133 7859 19136 7917
rect 19086 7856 19136 7859
rect 19150 31656 19200 31659
rect 19150 31598 19153 31656
rect 19197 31598 19200 31656
rect 760 6449 763 6507
rect 807 6449 810 6507
rect 760 6446 810 6449
rect 19150 6507 19200 31598
rect 19150 6449 19153 6507
rect 19197 6449 19200 6507
rect 19150 6446 19200 6449
rect 19214 31592 19264 31595
rect 19214 31534 19217 31592
rect 19261 31534 19264 31592
rect 696 6359 699 6417
rect 743 6359 746 6417
rect 696 6356 746 6359
rect 19214 6417 19264 31534
rect 19214 6359 19217 6417
rect 19261 6359 19264 6417
rect 19214 6356 19264 6359
rect 19278 31256 19328 31259
rect 19278 31198 19281 31256
rect 19325 31198 19328 31256
rect 12868 6201 12968 6204
rect 12868 6107 12871 6201
rect 12965 6107 12968 6201
rect 12868 5577 12968 6107
rect 12868 5483 12871 5577
rect 12965 5483 12968 5577
rect 12868 5480 12968 5483
rect 13006 6033 13106 6036
rect 13006 5939 13009 6033
rect 13103 5939 13106 6033
rect 13006 5577 13106 5939
rect 13006 5483 13009 5577
rect 13103 5483 13106 5577
rect 13006 5480 13106 5483
rect 13144 5865 13244 5868
rect 13144 5771 13147 5865
rect 13241 5771 13244 5865
rect 13144 5577 13244 5771
rect 13144 5483 13147 5577
rect 13241 5483 13244 5577
rect 13144 5480 13244 5483
rect 13282 5697 13382 5700
rect 13282 5603 13285 5697
rect 13379 5603 13382 5697
rect 13282 5577 13382 5603
rect 13282 5483 13285 5577
rect 13379 5483 13382 5577
rect 13282 5480 13382 5483
rect 632 4949 635 5007
rect 679 4949 682 5007
rect 632 4946 682 4949
rect 19278 5007 19328 31198
rect 19278 4949 19281 5007
rect 19325 4949 19328 5007
rect 19278 4946 19328 4949
rect 19342 31192 19392 31195
rect 19342 31134 19345 31192
rect 19389 31134 19392 31192
rect 568 4859 571 4917
rect 615 4859 618 4917
rect 568 4856 618 4859
rect 19342 4917 19392 31134
rect 19342 4859 19345 4917
rect 19389 4859 19392 4917
rect 19342 4856 19392 4859
rect 19406 30856 19456 30859
rect 19406 30798 19409 30856
rect 19453 30798 19456 30856
rect 504 3449 507 3507
rect 551 3449 554 3507
rect 504 3446 554 3449
rect 19406 3507 19456 30798
rect 19406 3449 19409 3507
rect 19453 3449 19456 3507
rect 19406 3446 19456 3449
rect 19470 30792 19520 30795
rect 19470 30734 19473 30792
rect 19517 30734 19520 30792
rect 440 3359 443 3417
rect 487 3359 490 3417
rect 440 3356 490 3359
rect 19470 3417 19520 30734
rect 19470 3359 19473 3417
rect 19517 3359 19520 3417
rect 19470 3356 19520 3359
rect 19534 30655 19584 30658
rect 19534 30597 19537 30655
rect 19581 30597 19584 30655
rect 376 1949 379 2007
rect 423 1949 426 2007
rect 376 1946 426 1949
rect 5903 2541 6000 2630
rect 5903 1980 5983 2541
rect 6083 2049 6400 2100
rect 6083 2023 6086 2049
rect 6138 2023 6400 2049
rect 6083 2020 6400 2023
rect 19534 2007 19584 30597
rect 5903 1977 12520 1980
rect 5903 1951 6814 1977
rect 6866 1951 7614 1977
rect 7666 1951 8414 1977
rect 8466 1951 9214 1977
rect 9266 1951 10014 1977
rect 10066 1951 10814 1977
rect 10866 1951 11614 1977
rect 11666 1951 12443 1977
rect 312 1859 315 1917
rect 359 1859 362 1917
rect 5903 1903 12443 1951
rect 12517 1903 12520 1977
rect 19534 1949 19537 2007
rect 19581 1949 19584 2007
rect 19534 1946 19584 1949
rect 19598 30591 19648 30594
rect 19598 30533 19601 30591
rect 19645 30533 19648 30591
rect 5903 1900 12520 1903
rect 19598 1917 19648 30533
rect 312 1856 362 1859
rect 6083 1870 6141 1873
rect 6083 1844 6086 1870
rect 6138 1844 6141 1870
rect 6373 1867 6396 1900
rect 6483 1870 6541 1873
rect 6083 1841 6141 1844
rect 6180 1854 6238 1857
rect 6180 1802 6183 1854
rect 6235 1802 6238 1854
rect 6483 1844 6486 1870
rect 6538 1844 6541 1870
rect 6773 1867 6796 1900
rect 6883 1870 6941 1873
rect 6483 1841 6541 1844
rect 6580 1854 6638 1857
rect 6180 1799 6238 1802
rect 6580 1802 6583 1854
rect 6635 1802 6638 1854
rect 6883 1844 6886 1870
rect 6938 1844 6941 1870
rect 7173 1867 7196 1900
rect 7283 1870 7341 1873
rect 6883 1841 6941 1844
rect 6980 1854 7038 1857
rect 6580 1799 6638 1802
rect 6980 1802 6983 1854
rect 7035 1802 7038 1854
rect 7283 1844 7286 1870
rect 7338 1844 7341 1870
rect 7573 1867 7596 1900
rect 7683 1870 7741 1873
rect 7283 1841 7341 1844
rect 7380 1854 7438 1857
rect 6980 1799 7038 1802
rect 7380 1802 7383 1854
rect 7435 1802 7438 1854
rect 7683 1844 7686 1870
rect 7738 1844 7741 1870
rect 7973 1867 7996 1900
rect 8083 1870 8141 1873
rect 7683 1841 7741 1844
rect 7780 1854 7838 1857
rect 7380 1799 7438 1802
rect 7780 1802 7783 1854
rect 7835 1802 7838 1854
rect 8083 1844 8086 1870
rect 8138 1844 8141 1870
rect 8373 1867 8396 1900
rect 8483 1870 8541 1873
rect 8083 1841 8141 1844
rect 8180 1854 8238 1857
rect 7780 1799 7838 1802
rect 8180 1802 8183 1854
rect 8235 1802 8238 1854
rect 8483 1844 8486 1870
rect 8538 1844 8541 1870
rect 8773 1867 8796 1900
rect 8883 1870 8941 1873
rect 8483 1841 8541 1844
rect 8580 1854 8638 1857
rect 8180 1799 8238 1802
rect 8580 1802 8583 1854
rect 8635 1802 8638 1854
rect 8883 1844 8886 1870
rect 8938 1844 8941 1870
rect 9173 1867 9196 1900
rect 9283 1870 9341 1873
rect 8883 1841 8941 1844
rect 8980 1854 9038 1857
rect 8580 1799 8638 1802
rect 8980 1802 8983 1854
rect 9035 1802 9038 1854
rect 9283 1844 9286 1870
rect 9338 1844 9341 1870
rect 9573 1867 9596 1900
rect 9683 1870 9741 1873
rect 9283 1841 9341 1844
rect 9380 1854 9438 1857
rect 8980 1799 9038 1802
rect 9380 1802 9383 1854
rect 9435 1802 9438 1854
rect 9683 1844 9686 1870
rect 9738 1844 9741 1870
rect 9973 1867 9996 1900
rect 10083 1870 10141 1873
rect 9683 1841 9741 1844
rect 9780 1854 9838 1857
rect 9380 1799 9438 1802
rect 9780 1802 9783 1854
rect 9835 1802 9838 1854
rect 10083 1844 10086 1870
rect 10138 1844 10141 1870
rect 10373 1867 10396 1900
rect 10483 1870 10541 1873
rect 10083 1841 10141 1844
rect 10180 1854 10238 1857
rect 9780 1799 9838 1802
rect 10180 1802 10183 1854
rect 10235 1802 10238 1854
rect 10483 1844 10486 1870
rect 10538 1844 10541 1870
rect 10773 1867 10796 1900
rect 10883 1870 10941 1873
rect 10483 1841 10541 1844
rect 10580 1854 10638 1857
rect 10180 1799 10238 1802
rect 10580 1802 10583 1854
rect 10635 1802 10638 1854
rect 10883 1844 10886 1870
rect 10938 1844 10941 1870
rect 11173 1867 11196 1900
rect 11283 1870 11341 1873
rect 10883 1841 10941 1844
rect 10980 1854 11038 1857
rect 10580 1799 10638 1802
rect 10980 1802 10983 1854
rect 11035 1802 11038 1854
rect 11283 1844 11286 1870
rect 11338 1844 11341 1870
rect 11573 1867 11596 1900
rect 11683 1870 11741 1873
rect 11283 1841 11341 1844
rect 11380 1854 11438 1857
rect 10980 1799 11038 1802
rect 11380 1802 11383 1854
rect 11435 1802 11438 1854
rect 11683 1844 11686 1870
rect 11738 1844 11741 1870
rect 11973 1867 11996 1900
rect 12083 1870 12141 1873
rect 11683 1841 11741 1844
rect 11780 1854 11838 1857
rect 11380 1799 11438 1802
rect 11780 1802 11783 1854
rect 11835 1802 11838 1854
rect 12083 1844 12086 1870
rect 12138 1844 12141 1870
rect 12373 1867 12396 1900
rect 19598 1859 19601 1917
rect 19645 1859 19648 1917
rect 12083 1841 12141 1844
rect 12180 1854 12238 1857
rect 19598 1856 19648 1859
rect 19662 30056 19712 30059
rect 19662 29998 19665 30056
rect 19709 29998 19712 30056
rect 11780 1799 11838 1802
rect 12180 1802 12183 1854
rect 12235 1802 12238 1854
rect 12180 1799 12238 1802
rect 6087 987 6116 990
rect 6087 593 6090 987
rect 6087 590 6116 593
rect 6487 987 6516 990
rect 6487 593 6490 987
rect 6487 590 6516 593
rect 6887 987 6916 990
rect 6887 593 6890 987
rect 6887 590 6916 593
rect 7287 987 7316 990
rect 7287 593 7290 987
rect 7287 590 7316 593
rect 7687 987 7716 990
rect 7687 593 7690 987
rect 7687 590 7716 593
rect 8087 987 8116 990
rect 8087 593 8090 987
rect 8087 590 8116 593
rect 8487 987 8516 990
rect 8487 593 8490 987
rect 8487 590 8516 593
rect 8887 987 8916 990
rect 8887 593 8890 987
rect 8887 590 8916 593
rect 9287 987 9316 990
rect 9287 593 9290 987
rect 9287 590 9316 593
rect 9687 987 9716 990
rect 9687 593 9690 987
rect 9687 590 9716 593
rect 10087 987 10116 990
rect 10087 593 10090 987
rect 10087 590 10116 593
rect 10487 987 10516 990
rect 10487 593 10490 987
rect 10487 590 10516 593
rect 10887 987 10916 990
rect 10887 593 10890 987
rect 10887 590 10916 593
rect 11287 987 11316 990
rect 11287 593 11290 987
rect 11287 590 11316 593
rect 11687 987 11716 990
rect 11687 593 11690 987
rect 11687 590 11716 593
rect 12087 987 12116 990
rect 12087 593 12090 987
rect 12087 590 12116 593
rect 248 449 251 507
rect 295 449 298 507
rect 248 446 298 449
rect 184 359 187 417
rect 231 359 234 417
rect 184 356 234 359
rect 1089 277 1139 280
rect 1089 233 1092 277
rect 1136 233 1139 277
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -220 -5 -140 0
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect -220 -80 -140 -75
rect 1027 -64 1059 -61
rect -18268 -984 -18236 -981
rect -18268 -1010 -18265 -984
rect -18239 -1010 -18236 -984
rect -18268 -1018 -18236 -1010
rect -18206 -1018 -18156 -80
rect -16268 -892 -16236 -889
rect -16268 -918 -16265 -892
rect -16239 -918 -16236 -892
rect -18014 -938 -17982 -935
rect -18014 -964 -18011 -938
rect -17985 -964 -17982 -938
rect -18014 -1018 -17982 -964
rect -16268 -1018 -16236 -918
rect -16206 -1018 -16156 -80
rect -14268 -800 -14236 -797
rect -14268 -826 -14265 -800
rect -14239 -826 -14236 -800
rect -16014 -846 -15982 -843
rect -16014 -872 -16011 -846
rect -15985 -872 -15982 -846
rect -16014 -1018 -15982 -872
rect -14268 -1018 -14236 -826
rect -14206 -1018 -14156 -80
rect -12268 -708 -12236 -705
rect -12268 -734 -12265 -708
rect -12239 -734 -12236 -708
rect -14014 -754 -13982 -751
rect -14014 -780 -14011 -754
rect -13985 -780 -13982 -754
rect -14014 -1018 -13982 -780
rect -12268 -1018 -12236 -734
rect -12206 -1018 -12156 -80
rect -10268 -616 -10236 -613
rect -10268 -642 -10265 -616
rect -10239 -642 -10236 -616
rect -12014 -662 -11982 -659
rect -12014 -688 -12011 -662
rect -11985 -688 -11982 -662
rect -12014 -1018 -11982 -688
rect -10268 -1018 -10236 -642
rect -10206 -1018 -10156 -80
rect -8268 -524 -8236 -521
rect -8268 -550 -8265 -524
rect -8239 -550 -8236 -524
rect -10014 -570 -9982 -567
rect -10014 -596 -10011 -570
rect -9985 -596 -9982 -570
rect -10014 -1018 -9982 -596
rect -8268 -1018 -8236 -550
rect -8206 -1018 -8156 -80
rect -6268 -432 -6236 -429
rect -6268 -458 -6265 -432
rect -6239 -458 -6236 -432
rect -8014 -478 -7982 -475
rect -8014 -504 -8011 -478
rect -7985 -504 -7982 -478
rect -8014 -1018 -7982 -504
rect -6268 -1018 -6236 -458
rect -6206 -1018 -6156 -80
rect -4268 -340 -4236 -337
rect -4268 -366 -4265 -340
rect -4239 -366 -4236 -340
rect -6014 -386 -5982 -383
rect -6014 -412 -6011 -386
rect -5985 -412 -5982 -386
rect -6014 -1018 -5982 -412
rect -4268 -1018 -4236 -366
rect -4206 -1018 -4156 -80
rect -2268 -248 -2236 -245
rect -2268 -274 -2265 -248
rect -2239 -274 -2236 -248
rect -4014 -294 -3982 -291
rect -4014 -320 -4011 -294
rect -3985 -320 -3982 -294
rect -4014 -1018 -3982 -320
rect -2268 -1018 -2236 -274
rect -2206 -1018 -2156 -80
rect -268 -156 -236 -153
rect -268 -182 -265 -156
rect -239 -182 -236 -156
rect -2014 -202 -1982 -199
rect -2014 -228 -2011 -202
rect -1985 -228 -1982 -202
rect -2014 -1018 -1982 -228
rect -268 -1018 -236 -182
rect -206 -1018 -156 -80
rect 1027 -90 1030 -64
rect 1056 -90 1059 -64
rect -14 -110 18 -107
rect -14 -136 -11 -110
rect 15 -136 18 -110
rect -14 -1018 18 -136
rect 1027 -1018 1059 -90
rect 1089 -1018 1139 233
rect 7281 166 7313 169
rect 7281 140 7284 166
rect 7310 140 7313 166
rect 7027 120 7059 123
rect 6281 74 6313 97
rect 6281 48 6284 74
rect 6310 48 6313 74
rect 6027 28 6059 31
rect 6027 2 6030 28
rect 6056 2 6059 28
rect 1281 -18 1313 -15
rect 1281 -44 1284 -18
rect 1310 -44 1313 -18
rect 1281 -1018 1313 -44
rect 6027 -1018 6059 2
rect 6281 -1018 6313 48
rect 7027 94 7030 120
rect 7056 94 7059 120
rect 7027 -1018 7059 94
rect 7281 -1018 7313 140
rect 7393 120 7425 557
rect 7447 166 7479 557
rect 7447 140 7450 166
rect 7476 140 7479 166
rect 7447 137 7479 140
rect 7393 94 7396 120
rect 7422 94 7425 120
rect 7393 91 7425 94
rect 7793 28 7825 557
rect 7847 74 7879 557
rect 7847 48 7850 74
rect 7876 48 7879 74
rect 7847 45 7879 48
rect 7793 2 7796 28
rect 7822 2 7825 28
rect 7793 -1 7825 2
rect 8193 -64 8225 557
rect 8247 -18 8279 557
rect 8247 -44 8250 -18
rect 8276 -44 8279 -18
rect 8247 -47 8279 -44
rect 8193 -90 8196 -64
rect 8222 -90 8225 -64
rect 8193 -93 8225 -90
rect 8593 -984 8625 557
rect 8647 -938 8679 557
rect 8993 -892 9025 557
rect 9047 -846 9079 557
rect 9393 -800 9425 557
rect 9447 -754 9479 557
rect 9793 -708 9825 557
rect 9847 -662 9879 557
rect 10193 -616 10225 557
rect 10247 -570 10279 557
rect 10593 -524 10625 557
rect 10647 -478 10679 557
rect 10993 -432 11025 557
rect 11047 -386 11079 557
rect 11393 -340 11425 557
rect 11447 -294 11479 557
rect 11793 -248 11825 557
rect 11847 -202 11879 557
rect 12193 -156 12225 557
rect 12247 -110 12279 557
rect 19662 507 19712 29998
rect 19662 449 19665 507
rect 19709 449 19712 507
rect 19662 446 19712 449
rect 19726 29992 19776 29995
rect 19726 29934 19729 29992
rect 19773 29934 19776 29992
rect 19726 417 19776 29934
rect 19726 359 19729 417
rect 19773 359 19776 417
rect 19726 356 19776 359
rect 20100 -5 20180 0
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
rect 12247 -136 12250 -110
rect 12276 -136 12279 -110
rect 12247 -139 12279 -136
rect 19941 -110 19973 -107
rect 19941 -136 19944 -110
rect 19970 -136 19973 -110
rect 12193 -182 12196 -156
rect 12222 -182 12225 -156
rect 12193 -185 12225 -182
rect 11847 -228 11850 -202
rect 11876 -228 11879 -202
rect 11847 -231 11879 -228
rect 11793 -274 11796 -248
rect 11822 -274 11825 -248
rect 11793 -277 11825 -274
rect 11447 -320 11450 -294
rect 11476 -320 11479 -294
rect 11447 -323 11479 -320
rect 11393 -366 11396 -340
rect 11422 -366 11425 -340
rect 11393 -369 11425 -366
rect 11047 -412 11050 -386
rect 11076 -412 11079 -386
rect 11047 -415 11079 -412
rect 10993 -458 10996 -432
rect 11022 -458 11025 -432
rect 10993 -461 11025 -458
rect 10647 -504 10650 -478
rect 10676 -504 10679 -478
rect 10647 -507 10679 -504
rect 10593 -550 10596 -524
rect 10622 -550 10625 -524
rect 10593 -553 10625 -550
rect 10247 -596 10250 -570
rect 10276 -596 10279 -570
rect 10247 -599 10279 -596
rect 10193 -642 10196 -616
rect 10222 -642 10225 -616
rect 10193 -645 10225 -642
rect 9847 -688 9850 -662
rect 9876 -688 9879 -662
rect 9847 -691 9879 -688
rect 9793 -734 9796 -708
rect 9822 -734 9825 -708
rect 9793 -737 9825 -734
rect 9447 -780 9450 -754
rect 9476 -780 9479 -754
rect 9447 -783 9479 -780
rect 9393 -826 9396 -800
rect 9422 -826 9425 -800
rect 9393 -829 9425 -826
rect 9047 -872 9050 -846
rect 9076 -872 9079 -846
rect 9047 -875 9079 -872
rect 8993 -918 8996 -892
rect 9022 -918 9025 -892
rect 8993 -921 9025 -918
rect 8647 -964 8650 -938
rect 8676 -964 8679 -938
rect 8647 -967 8679 -964
rect 8593 -1010 8596 -984
rect 8622 -1010 8625 -984
rect 8593 -1013 8625 -1010
rect 19941 -1018 19973 -136
rect 20115 -1018 20165 -80
rect 20195 -156 20227 -153
rect 20195 -182 20198 -156
rect 20224 -182 20227 -156
rect 20195 -1018 20227 -182
rect 21941 -202 21973 -199
rect 21941 -228 21944 -202
rect 21970 -228 21973 -202
rect 21941 -1018 21973 -228
rect 22115 -1018 22165 -80
rect 22195 -248 22227 -245
rect 22195 -274 22198 -248
rect 22224 -274 22227 -248
rect 22195 -1018 22227 -274
rect 23941 -294 23973 -291
rect 23941 -320 23944 -294
rect 23970 -320 23973 -294
rect 23941 -1018 23973 -320
rect 24115 -1018 24165 -80
rect 24195 -340 24227 -337
rect 24195 -366 24198 -340
rect 24224 -366 24227 -340
rect 24195 -1018 24227 -366
rect 25941 -386 25973 -383
rect 25941 -412 25944 -386
rect 25970 -412 25973 -386
rect 25941 -1018 25973 -412
rect 26115 -1018 26165 -80
rect 26195 -432 26227 -429
rect 26195 -458 26198 -432
rect 26224 -458 26227 -432
rect 26195 -1018 26227 -458
rect 27941 -478 27973 -475
rect 27941 -504 27944 -478
rect 27970 -504 27973 -478
rect 27941 -1018 27973 -504
rect 28115 -1018 28165 -80
rect 28195 -524 28227 -521
rect 28195 -550 28198 -524
rect 28224 -550 28227 -524
rect 28195 -1018 28227 -550
rect 29941 -570 29973 -567
rect 29941 -596 29944 -570
rect 29970 -596 29973 -570
rect 29941 -1018 29973 -596
rect 30115 -1018 30165 -80
rect 30195 -616 30227 -613
rect 30195 -642 30198 -616
rect 30224 -642 30227 -616
rect 30195 -1018 30227 -642
rect 31941 -662 31973 -659
rect 31941 -688 31944 -662
rect 31970 -688 31973 -662
rect 31941 -1018 31973 -688
rect 32115 -1018 32165 -80
rect 32195 -708 32227 -705
rect 32195 -734 32198 -708
rect 32224 -734 32227 -708
rect 32195 -1018 32227 -734
rect 33941 -754 33973 -751
rect 33941 -780 33944 -754
rect 33970 -780 33973 -754
rect 33941 -1018 33973 -780
rect 34115 -1018 34165 -80
rect 34195 -800 34227 -797
rect 34195 -826 34198 -800
rect 34224 -826 34227 -800
rect 34195 -1018 34227 -826
rect 35941 -846 35973 -843
rect 35941 -872 35944 -846
rect 35970 -872 35973 -846
rect 35941 -1018 35973 -872
rect 36115 -1018 36165 -80
rect 36195 -892 36227 -889
rect 36195 -918 36198 -892
rect 36224 -918 36227 -892
rect 36195 -1018 36227 -918
rect 37941 -938 37973 -935
rect 37941 -964 37944 -938
rect 37970 -964 37973 -938
rect 37941 -1018 37973 -964
rect 38115 -1018 38165 -80
rect 38195 -984 38227 -981
rect 38195 -1010 38198 -984
rect 38224 -1010 38227 -984
rect 38195 -1018 38227 -1010
rect -17943 -1100 -17817 -1097
rect -17943 -1220 -17940 -1100
rect -17820 -1220 -17817 -1100
rect -17943 -1223 -17817 -1220
rect -15943 -1100 -15817 -1097
rect -15943 -1220 -15940 -1100
rect -15820 -1220 -15817 -1100
rect -15943 -1223 -15817 -1220
rect -13943 -1100 -13817 -1097
rect -13943 -1220 -13940 -1100
rect -13820 -1220 -13817 -1100
rect -13943 -1223 -13817 -1220
rect -11943 -1100 -11817 -1097
rect -11943 -1220 -11940 -1100
rect -11820 -1220 -11817 -1100
rect -11943 -1223 -11817 -1220
rect -9943 -1100 -9817 -1097
rect -9943 -1220 -9940 -1100
rect -9820 -1220 -9817 -1100
rect -9943 -1223 -9817 -1220
rect -7943 -1100 -7817 -1097
rect -7943 -1220 -7940 -1100
rect -7820 -1220 -7817 -1100
rect -7943 -1223 -7817 -1220
rect -5943 -1100 -5817 -1097
rect -5943 -1220 -5940 -1100
rect -5820 -1220 -5817 -1100
rect -5943 -1223 -5817 -1220
rect -3943 -1100 -3817 -1097
rect -3943 -1220 -3940 -1100
rect -3820 -1220 -3817 -1100
rect -3943 -1223 -3817 -1220
rect -1943 -1100 -1817 -1097
rect -1943 -1220 -1940 -1100
rect -1820 -1220 -1817 -1100
rect -1943 -1223 -1817 -1220
rect 57 -1100 183 -1097
rect 57 -1220 60 -1100
rect 180 -1220 183 -1100
rect 57 -1223 183 -1220
rect 1352 -1100 1478 -1097
rect 1352 -1220 1355 -1100
rect 1475 -1220 1478 -1100
rect 1352 -1223 1478 -1220
rect 6352 -1100 6478 -1097
rect 6352 -1220 6355 -1100
rect 6475 -1220 6478 -1100
rect 6352 -1223 6478 -1220
rect 7352 -1100 7478 -1097
rect 7352 -1220 7355 -1100
rect 7475 -1220 7478 -1100
rect 7352 -1223 7478 -1220
rect 19773 -1100 19899 -1097
rect 19773 -1220 19776 -1100
rect 19896 -1220 19899 -1100
rect 19773 -1223 19899 -1220
rect 21773 -1100 21899 -1097
rect 21773 -1220 21776 -1100
rect 21896 -1220 21899 -1100
rect 21773 -1223 21899 -1220
rect 23773 -1100 23899 -1097
rect 23773 -1220 23776 -1100
rect 23896 -1220 23899 -1100
rect 23773 -1223 23899 -1220
rect 25773 -1100 25899 -1097
rect 25773 -1220 25776 -1100
rect 25896 -1220 25899 -1100
rect 25773 -1223 25899 -1220
rect 27773 -1100 27899 -1097
rect 27773 -1220 27776 -1100
rect 27896 -1220 27899 -1100
rect 27773 -1223 27899 -1220
rect 29773 -1100 29899 -1097
rect 29773 -1220 29776 -1100
rect 29896 -1220 29899 -1100
rect 29773 -1223 29899 -1220
rect 31773 -1100 31899 -1097
rect 31773 -1220 31776 -1100
rect 31896 -1220 31899 -1100
rect 31773 -1223 31899 -1220
rect 33773 -1100 33899 -1097
rect 33773 -1220 33776 -1100
rect 33896 -1220 33899 -1100
rect 33773 -1223 33899 -1220
rect 35773 -1100 35899 -1097
rect 35773 -1220 35776 -1100
rect 35896 -1220 35899 -1100
rect 35773 -1223 35899 -1220
rect 37773 -1100 37899 -1097
rect 37773 -1220 37776 -1100
rect 37896 -1220 37899 -1100
rect 37773 -1223 37899 -1220
rect -18443 -1710 -18313 -1705
rect -18443 -1830 -18438 -1710
rect -18318 -1830 -18313 -1710
rect -16443 -1710 -16313 -1705
rect -18443 -1835 -18313 -1830
rect -18090 -2000 -18030 -1720
rect -16443 -1830 -16438 -1710
rect -16318 -1830 -16313 -1710
rect -14443 -1710 -14313 -1705
rect -16443 -1835 -16313 -1830
rect -16090 -2000 -16030 -1720
rect -14443 -1830 -14438 -1710
rect -14318 -1830 -14313 -1710
rect -12443 -1710 -12313 -1705
rect -14443 -1835 -14313 -1830
rect -14090 -2000 -14030 -1720
rect -12443 -1830 -12438 -1710
rect -12318 -1830 -12313 -1710
rect -10443 -1710 -10313 -1705
rect -12443 -1835 -12313 -1830
rect -12090 -2000 -12030 -1720
rect -10443 -1830 -10438 -1710
rect -10318 -1830 -10313 -1710
rect -8443 -1710 -8313 -1705
rect -10443 -1835 -10313 -1830
rect -10090 -2000 -10030 -1720
rect -8443 -1830 -8438 -1710
rect -8318 -1830 -8313 -1710
rect -6443 -1710 -6313 -1705
rect -8443 -1835 -8313 -1830
rect -8090 -2000 -8030 -1720
rect -6443 -1830 -6438 -1710
rect -6318 -1830 -6313 -1710
rect -4443 -1710 -4313 -1705
rect -6443 -1835 -6313 -1830
rect -6090 -2000 -6030 -1720
rect -4443 -1830 -4438 -1710
rect -4318 -1830 -4313 -1710
rect -2443 -1710 -2313 -1705
rect -4443 -1835 -4313 -1830
rect -4090 -2000 -4030 -1720
rect -2443 -1830 -2438 -1710
rect -2318 -1830 -2313 -1710
rect -443 -1710 -313 -1705
rect -2443 -1835 -2313 -1830
rect -2090 -2000 -2030 -1720
rect -443 -1830 -438 -1710
rect -318 -1830 -313 -1710
rect 852 -1710 982 -1705
rect -443 -1835 -313 -1830
rect -90 -2000 -30 -1720
rect 852 -1830 857 -1710
rect 977 -1830 982 -1710
rect 5852 -1710 5982 -1705
rect 852 -1835 982 -1830
rect 1205 -2000 1265 -1720
rect 5852 -1830 5857 -1710
rect 5977 -1770 5982 -1710
rect 6089 -1770 6139 -1697
rect 6852 -1710 6982 -1705
rect 5977 -1830 6139 -1770
rect 5852 -1835 6139 -1830
rect 6205 -2000 6265 -1720
rect 6852 -1830 6857 -1710
rect 6977 -1830 6982 -1710
rect 20255 -1710 20385 -1705
rect 6852 -1835 6982 -1830
rect 7205 -2000 7265 -1720
rect 19990 -2000 20050 -1730
rect 20255 -1830 20260 -1710
rect 20380 -1830 20385 -1710
rect 22255 -1710 22385 -1705
rect 20255 -1835 20385 -1830
rect 21990 -2000 22050 -1730
rect 22255 -1830 22260 -1710
rect 22380 -1830 22385 -1710
rect 24255 -1710 24385 -1705
rect 22255 -1835 22385 -1830
rect 23990 -2000 24050 -1730
rect 24255 -1830 24260 -1710
rect 24380 -1830 24385 -1710
rect 26255 -1710 26385 -1705
rect 24255 -1835 24385 -1830
rect 25990 -2000 26050 -1730
rect 26255 -1830 26260 -1710
rect 26380 -1830 26385 -1710
rect 28255 -1710 28385 -1705
rect 26255 -1835 26385 -1830
rect 27990 -2000 28050 -1730
rect 28255 -1830 28260 -1710
rect 28380 -1830 28385 -1710
rect 30255 -1710 30385 -1705
rect 28255 -1835 28385 -1830
rect 29990 -2000 30050 -1730
rect 30255 -1830 30260 -1710
rect 30380 -1830 30385 -1710
rect 32255 -1710 32385 -1705
rect 30255 -1835 30385 -1830
rect 31990 -2000 32050 -1730
rect 32255 -1830 32260 -1710
rect 32380 -1830 32385 -1710
rect 34255 -1710 34385 -1705
rect 32255 -1835 32385 -1830
rect 33990 -2000 34050 -1730
rect 34255 -1830 34260 -1710
rect 34380 -1830 34385 -1710
rect 36255 -1710 36385 -1705
rect 34255 -1835 34385 -1830
rect 35990 -2000 36050 -1730
rect 36255 -1830 36260 -1710
rect 36380 -1830 36385 -1710
rect 38255 -1710 38385 -1705
rect 36255 -1835 36385 -1830
rect 37990 -2000 38050 -1730
rect 38255 -1830 38260 -1710
rect 38380 -1830 38385 -1710
rect 38255 -1835 38385 -1830
rect -18090 -2010 7390 -2000
rect -18090 -2190 4410 -2010
rect 4790 -2190 7390 -2010
rect -18090 -2200 7390 -2190
rect 17200 -2020 38050 -2000
rect 17200 -2180 17220 -2020
rect 17780 -2180 38050 -2020
rect 17200 -2200 38050 -2180
<< via1 >>
rect 3259 43963 3303 44021
rect 16657 43963 16701 44021
rect 3259 41584 3303 41642
rect 3323 43873 3367 43931
rect 16593 43873 16637 43931
rect 3323 41520 3367 41578
rect 3387 42463 3431 42521
rect 16529 42463 16573 42521
rect 3387 41184 3431 41242
rect 3451 42373 3495 42431
rect 16465 42373 16509 42431
rect 5090 41793 5170 41871
rect 14790 41793 14870 41871
rect 3680 41598 3724 41642
rect 3680 41534 3724 41578
rect 4992 41535 5044 41587
rect 3853 41447 4257 41473
rect 5034 41438 5060 41496
rect 5213 41438 5239 41496
rect 14721 41438 14747 41496
rect 3680 41198 3724 41242
rect 3451 41120 3495 41178
rect 3680 41134 3724 41178
rect 4992 41135 5044 41187
rect 3853 41047 4257 41073
rect 5034 41038 5060 41096
rect 3515 40963 3559 41021
rect 16236 41598 16280 41642
rect 14916 41535 14968 41587
rect 16236 41534 16280 41578
rect 14900 41438 14926 41496
rect 15703 41447 16107 41473
rect 5213 41038 5239 41096
rect 14721 41038 14747 41096
rect 16236 41198 16280 41242
rect 14916 41135 14968 41187
rect 16236 41134 16280 41178
rect 16657 41584 16701 41642
rect 16593 41520 16637 41578
rect 16529 41184 16573 41242
rect 16465 41120 16509 41178
rect 14900 41038 14926 41096
rect 15703 41047 16107 41073
rect 5141 40960 5167 41018
rect 5320 40960 5346 41018
rect 14614 40960 14640 41018
rect 14793 40960 14819 41018
rect 3515 40784 3559 40842
rect 3579 40873 3623 40931
rect 3680 40798 3724 40842
rect 3579 40720 3623 40778
rect 3680 40734 3724 40778
rect 4992 40735 5044 40787
rect 3853 40647 4257 40673
rect 5034 40638 5060 40696
rect 16401 40963 16445 41021
rect 5213 40638 5239 40696
rect 14721 40638 14747 40696
rect 3579 40398 3623 40456
rect 3515 40334 3559 40392
rect 3451 39998 3495 40056
rect 3387 39934 3431 39992
rect 3323 39598 3367 39656
rect 3259 39534 3303 39592
rect 3195 39198 3239 39256
rect 3131 39134 3175 39192
rect 3067 38798 3111 38856
rect 3003 38734 3047 38792
rect 2939 38398 2983 38456
rect 2875 38334 2919 38392
rect 2811 38097 2855 38155
rect 2747 38033 2791 38091
rect 2683 37598 2727 37656
rect 2619 37534 2663 37592
rect 2555 37198 2599 37256
rect 2491 37134 2535 37192
rect 2427 36798 2471 36856
rect 2363 36734 2407 36792
rect 2299 36597 2343 36655
rect 2235 36533 2279 36591
rect 2171 35998 2215 36056
rect 2107 35934 2151 35992
rect 2043 35598 2087 35656
rect 1979 35534 2023 35592
rect 1915 35198 1959 35256
rect 1851 35134 1895 35192
rect 1787 34795 1831 34853
rect 1723 34731 1767 34789
rect 1659 34398 1703 34456
rect 1595 34334 1639 34392
rect 1531 33998 1575 34056
rect 1467 33934 1511 33992
rect 1403 33598 1447 33656
rect 1339 33534 1383 33592
rect 1275 33198 1319 33256
rect 1211 33134 1255 33192
rect 1147 32798 1191 32856
rect 1083 32734 1127 32792
rect 1019 32398 1063 32456
rect 955 32334 999 32392
rect 891 32091 935 32149
rect 827 32027 871 32085
rect 763 31598 807 31656
rect 699 31534 743 31592
rect 635 31198 679 31256
rect 571 31134 615 31192
rect 507 30798 551 30856
rect 443 30734 487 30792
rect 379 30597 423 30655
rect 315 30533 359 30591
rect 251 29998 295 30056
rect 187 29934 231 29992
rect 3680 40398 3724 40442
rect 3680 40334 3724 40378
rect 4992 40335 5044 40387
rect 3853 40247 4257 40273
rect 5034 40238 5060 40296
rect 16337 40873 16381 40931
rect 16236 40798 16280 40842
rect 14916 40735 14968 40787
rect 16236 40734 16280 40778
rect 16401 40784 16445 40842
rect 16337 40720 16381 40778
rect 14900 40638 14926 40696
rect 15703 40647 16107 40673
rect 5213 40238 5239 40296
rect 14721 40238 14747 40296
rect 16236 40398 16280 40442
rect 16337 40398 16381 40456
rect 14916 40335 14968 40387
rect 16236 40334 16280 40378
rect 14900 40238 14926 40296
rect 15703 40247 16107 40273
rect 5141 40160 5167 40218
rect 5320 40160 5346 40218
rect 14614 40160 14640 40218
rect 14793 40160 14819 40218
rect 3680 39998 3724 40042
rect 3680 39934 3724 39978
rect 4992 39935 5044 39987
rect 3853 39847 4257 39873
rect 5034 39838 5060 39896
rect 5213 39838 5239 39896
rect 14721 39838 14747 39896
rect 3680 39598 3724 39642
rect 3680 39534 3724 39578
rect 4992 39535 5044 39587
rect 3579 39449 3623 39507
rect 3853 39447 4257 39473
rect 5034 39438 5060 39496
rect 3515 39359 3559 39417
rect 16236 39998 16280 40042
rect 14916 39935 14968 39987
rect 16236 39934 16280 39978
rect 14900 39838 14926 39896
rect 15703 39847 16107 39873
rect 5213 39438 5239 39496
rect 14721 39438 14747 39496
rect 16236 39598 16280 39642
rect 14916 39535 14968 39587
rect 16236 39534 16280 39578
rect 14900 39438 14926 39496
rect 15703 39447 16107 39473
rect 16337 39449 16381 39507
rect 16401 40334 16445 40392
rect 5141 39360 5167 39418
rect 5320 39360 5346 39418
rect 14614 39360 14640 39418
rect 14793 39360 14819 39418
rect 3680 39198 3724 39242
rect 3680 39134 3724 39178
rect 4992 39135 5044 39187
rect 3853 39047 4257 39073
rect 5034 39038 5060 39096
rect 16401 39359 16445 39417
rect 16465 39998 16509 40056
rect 5213 39038 5239 39096
rect 14721 39038 14747 39096
rect 3680 38798 3724 38842
rect 3680 38734 3724 38778
rect 4992 38735 5044 38787
rect 3853 38647 4257 38673
rect 5034 38638 5060 38696
rect 16236 39198 16280 39242
rect 14916 39135 14968 39187
rect 16236 39134 16280 39178
rect 14900 39038 14926 39096
rect 15703 39047 16107 39073
rect 5213 38638 5239 38696
rect 14721 38638 14747 38696
rect 16236 38798 16280 38842
rect 14916 38735 14968 38787
rect 16236 38734 16280 38778
rect 14900 38638 14926 38696
rect 15703 38647 16107 38673
rect 5141 38560 5167 38618
rect 5320 38560 5346 38618
rect 14614 38560 14640 38618
rect 14793 38560 14819 38618
rect 3680 38398 3724 38442
rect 3680 38334 3724 38378
rect 4992 38335 5044 38387
rect 3853 38247 4257 38273
rect 5034 38238 5060 38296
rect 5213 38238 5239 38296
rect 14721 38238 14747 38296
rect 3451 37949 3495 38007
rect 3680 37998 3724 38042
rect 3680 37934 3724 37978
rect 4992 37935 5044 37987
rect 3387 37859 3431 37917
rect 3853 37847 4257 37873
rect 5034 37838 5060 37896
rect 16236 38398 16280 38442
rect 14916 38335 14968 38387
rect 16236 38334 16280 38378
rect 14900 38238 14926 38296
rect 15703 38247 16107 38273
rect 5213 37838 5239 37896
rect 14721 37838 14747 37896
rect 16236 37998 16280 38042
rect 14916 37935 14968 37987
rect 16236 37934 16280 37978
rect 16465 37949 16509 38007
rect 16529 39934 16573 39992
rect 14900 37838 14926 37896
rect 15703 37847 16107 37873
rect 16529 37859 16573 37917
rect 16593 39598 16637 39656
rect 5141 37760 5167 37818
rect 5320 37760 5346 37818
rect 14614 37760 14640 37818
rect 14793 37760 14819 37818
rect 3680 37598 3724 37642
rect 3680 37534 3724 37578
rect 4992 37535 5044 37587
rect 3853 37447 4257 37473
rect 5034 37438 5060 37496
rect 5213 37438 5239 37496
rect 14721 37438 14747 37496
rect 3680 37198 3724 37242
rect 3680 37134 3724 37178
rect 4992 37135 5044 37187
rect 3853 37047 4257 37073
rect 5034 37038 5060 37096
rect 16236 37598 16280 37642
rect 14916 37535 14968 37587
rect 16236 37534 16280 37578
rect 14900 37438 14926 37496
rect 15703 37447 16107 37473
rect 5213 37038 5239 37096
rect 14721 37038 14747 37096
rect 16236 37198 16280 37242
rect 14916 37135 14968 37187
rect 16236 37134 16280 37178
rect 14900 37038 14926 37096
rect 15703 37047 16107 37073
rect 5141 36960 5167 37018
rect 5320 36960 5346 37018
rect 14614 36960 14640 37018
rect 14793 36960 14819 37018
rect 3680 36798 3724 36842
rect 3680 36734 3724 36778
rect 4992 36735 5044 36787
rect 3853 36647 4257 36673
rect 5034 36638 5060 36696
rect 5213 36638 5239 36696
rect 14721 36638 14747 36696
rect 3323 36449 3367 36507
rect 3259 36359 3303 36417
rect 3680 36398 3724 36442
rect 3680 36334 3724 36378
rect 4992 36335 5044 36387
rect 3853 36247 4257 36273
rect 5034 36238 5060 36296
rect 16236 36798 16280 36842
rect 14916 36735 14968 36787
rect 16236 36734 16280 36778
rect 14900 36638 14926 36696
rect 15703 36647 16107 36673
rect 5213 36238 5239 36296
rect 14721 36238 14747 36296
rect 16593 36449 16637 36507
rect 16657 39534 16701 39592
rect 16236 36398 16280 36442
rect 14916 36335 14968 36387
rect 16236 36334 16280 36378
rect 16657 36359 16701 36417
rect 16721 39198 16765 39256
rect 14900 36238 14926 36296
rect 15703 36247 16107 36273
rect 5141 36160 5167 36218
rect 5320 36160 5346 36218
rect 14614 36160 14640 36218
rect 14793 36160 14819 36218
rect 3680 35998 3724 36042
rect 3680 35934 3724 35978
rect 4992 35935 5044 35987
rect 3853 35847 4257 35873
rect 5034 35838 5060 35896
rect 5213 35838 5239 35896
rect 14721 35838 14747 35896
rect 3680 35598 3724 35642
rect 3680 35534 3724 35578
rect 4992 35535 5044 35587
rect 3853 35447 4257 35473
rect 5034 35438 5060 35496
rect 16236 35998 16280 36042
rect 14916 35935 14968 35987
rect 16236 35934 16280 35978
rect 14900 35838 14926 35896
rect 15703 35847 16107 35873
rect 5213 35438 5239 35496
rect 14721 35438 14747 35496
rect 16236 35598 16280 35642
rect 14916 35535 14968 35587
rect 16236 35534 16280 35578
rect 14900 35438 14926 35496
rect 15703 35447 16107 35473
rect 5141 35360 5167 35418
rect 5320 35360 5346 35418
rect 14614 35360 14640 35418
rect 14793 35360 14819 35418
rect 3680 35198 3724 35242
rect 3680 35134 3724 35178
rect 4992 35135 5044 35187
rect 3853 35047 4257 35073
rect 5034 35038 5060 35096
rect 3195 34949 3239 35007
rect 5213 35038 5239 35096
rect 14721 35038 14747 35096
rect 3131 34859 3175 34917
rect 3680 34798 3724 34842
rect 3680 34734 3724 34778
rect 4992 34735 5044 34787
rect 3853 34647 4257 34673
rect 5034 34638 5060 34696
rect 16236 35198 16280 35242
rect 14916 35135 14968 35187
rect 16236 35134 16280 35178
rect 14900 35038 14926 35096
rect 15703 35047 16107 35073
rect 16721 34949 16765 35007
rect 16785 39134 16829 39192
rect 5213 34638 5239 34696
rect 14721 34638 14747 34696
rect 16785 34859 16829 34917
rect 16849 38798 16893 38856
rect 16236 34798 16280 34842
rect 14916 34735 14968 34787
rect 16236 34734 16280 34778
rect 14900 34638 14926 34696
rect 15703 34647 16107 34673
rect 5141 34560 5167 34618
rect 5320 34560 5346 34618
rect 14614 34560 14640 34618
rect 14793 34560 14819 34618
rect 3680 34398 3724 34442
rect 3680 34334 3724 34378
rect 4992 34335 5044 34387
rect 3853 34247 4257 34273
rect 5034 34238 5060 34296
rect 5213 34238 5239 34296
rect 14721 34238 14747 34296
rect 3680 33998 3724 34042
rect 3680 33934 3724 33978
rect 4992 33935 5044 33987
rect 3853 33847 4257 33873
rect 5034 33838 5060 33896
rect 16236 34398 16280 34442
rect 14916 34335 14968 34387
rect 16236 34334 16280 34378
rect 14900 34238 14926 34296
rect 15703 34247 16107 34273
rect 5213 33838 5239 33896
rect 14721 33838 14747 33896
rect 16236 33998 16280 34042
rect 14916 33935 14968 33987
rect 16236 33934 16280 33978
rect 14900 33838 14926 33896
rect 15703 33847 16107 33873
rect 5141 33760 5167 33818
rect 5320 33760 5346 33818
rect 14614 33760 14640 33818
rect 14793 33760 14819 33818
rect 3680 33598 3724 33642
rect 3680 33534 3724 33578
rect 4992 33535 5044 33587
rect 3067 33449 3111 33507
rect 3853 33447 4257 33473
rect 5034 33438 5060 33496
rect 3003 33359 3047 33417
rect 5213 33438 5239 33496
rect 14721 33438 14747 33496
rect 3680 33198 3724 33242
rect 3680 33134 3724 33178
rect 4992 33135 5044 33187
rect 3853 33047 4257 33073
rect 5034 33038 5060 33096
rect 16236 33598 16280 33642
rect 14916 33535 14968 33587
rect 16236 33534 16280 33578
rect 14900 33438 14926 33496
rect 15703 33447 16107 33473
rect 16849 33449 16893 33507
rect 16913 38734 16957 38792
rect 16913 33359 16957 33417
rect 16977 38398 17021 38456
rect 5213 33038 5239 33096
rect 14721 33038 14747 33096
rect 16236 33198 16280 33242
rect 14916 33135 14968 33187
rect 16236 33134 16280 33178
rect 14900 33038 14926 33096
rect 15703 33047 16107 33073
rect 5141 32960 5167 33018
rect 5320 32960 5346 33018
rect 14614 32960 14640 33018
rect 14793 32960 14819 33018
rect 3680 32798 3724 32842
rect 3680 32734 3724 32778
rect 4992 32735 5044 32787
rect 3853 32647 4257 32673
rect 5034 32638 5060 32696
rect 5213 32638 5239 32696
rect 14721 32638 14747 32696
rect 3680 32398 3724 32442
rect 3680 32334 3724 32378
rect 4992 32335 5044 32387
rect 3853 32247 4257 32273
rect 5034 32238 5060 32296
rect 16236 32798 16280 32842
rect 14916 32735 14968 32787
rect 16236 32734 16280 32778
rect 14900 32638 14926 32696
rect 15703 32647 16107 32673
rect 5213 32238 5239 32296
rect 14721 32238 14747 32296
rect 16236 32398 16280 32442
rect 14916 32335 14968 32387
rect 16236 32334 16280 32378
rect 14900 32238 14926 32296
rect 15703 32247 16107 32273
rect 5141 32160 5167 32218
rect 5320 32160 5346 32218
rect 14614 32160 14640 32218
rect 14793 32160 14819 32218
rect 2939 31949 2983 32007
rect 3680 31998 3724 32042
rect 3680 31934 3724 31978
rect 4992 31935 5044 31987
rect 2875 31859 2919 31917
rect 3853 31847 4257 31873
rect 5034 31838 5060 31896
rect 5213 31838 5239 31896
rect 14721 31838 14747 31896
rect 3680 31598 3724 31642
rect 3680 31534 3724 31578
rect 4992 31535 5044 31587
rect 3853 31447 4257 31473
rect 5034 31438 5060 31496
rect 16236 31998 16280 32042
rect 14916 31935 14968 31987
rect 16236 31934 16280 31978
rect 16977 31949 17021 32007
rect 17041 38334 17085 38392
rect 14900 31838 14926 31896
rect 15703 31847 16107 31873
rect 17041 31859 17085 31917
rect 17105 38097 17149 38155
rect 5213 31438 5239 31496
rect 14721 31438 14747 31496
rect 16236 31598 16280 31642
rect 14916 31535 14968 31587
rect 16236 31534 16280 31578
rect 14900 31438 14926 31496
rect 15703 31447 16107 31473
rect 5141 31360 5167 31418
rect 5320 31360 5346 31418
rect 14614 31360 14640 31418
rect 14793 31360 14819 31418
rect 3680 31198 3724 31242
rect 3680 31134 3724 31178
rect 4992 31135 5044 31187
rect 3853 31047 4257 31073
rect 5034 31038 5060 31096
rect 5213 31038 5239 31096
rect 14721 31038 14747 31096
rect 3680 30798 3724 30842
rect 3680 30734 3724 30778
rect 4992 30735 5044 30787
rect 3853 30647 4257 30673
rect 5034 30638 5060 30696
rect 16236 31198 16280 31242
rect 14916 31135 14968 31187
rect 16236 31134 16280 31178
rect 14900 31038 14926 31096
rect 15703 31047 16107 31073
rect 5213 30638 5239 30696
rect 14721 30638 14747 30696
rect 16236 30798 16280 30842
rect 14916 30735 14968 30787
rect 16236 30734 16280 30778
rect 14900 30638 14926 30696
rect 15703 30647 16107 30673
rect 5141 30560 5167 30618
rect 5320 30560 5346 30618
rect 14614 30560 14640 30618
rect 14793 30560 14819 30618
rect 2811 30449 2855 30507
rect 2747 30359 2791 30417
rect 3680 30398 3724 30442
rect 3680 30334 3724 30378
rect 4992 30335 5044 30387
rect 3853 30247 4257 30273
rect 5034 30238 5060 30296
rect 5213 30238 5239 30296
rect 14721 30238 14747 30296
rect 3680 29998 3724 30042
rect 3680 29934 3724 29978
rect 4992 29935 5044 29987
rect 3853 29847 4257 29873
rect 5034 29838 5060 29896
rect 17105 30449 17149 30507
rect 17169 38033 17213 38091
rect 16236 30398 16280 30442
rect 14916 30335 14968 30387
rect 16236 30334 16280 30378
rect 17169 30359 17213 30417
rect 17233 37598 17277 37656
rect 14900 30238 14926 30296
rect 15703 30247 16107 30273
rect 5213 29838 5239 29896
rect 14721 29838 14747 29896
rect 16236 29998 16280 30042
rect 14916 29935 14968 29987
rect 16236 29934 16280 29978
rect 14900 29838 14926 29896
rect 15703 29847 16107 29873
rect 5141 29760 5167 29818
rect 5320 29760 5346 29818
rect 14614 29760 14640 29818
rect 14793 29760 14819 29818
rect 3680 29598 3724 29642
rect 3680 29534 3724 29578
rect 4992 29535 5044 29587
rect 3853 29447 4257 29473
rect 5034 29438 5060 29496
rect 5213 29438 5239 29496
rect 14721 29438 14747 29496
rect 16236 29598 16280 29642
rect 14916 29535 14968 29587
rect 16236 29534 16280 29578
rect 14900 29438 14926 29496
rect 15703 29447 16107 29473
rect 3680 29198 3724 29242
rect 3680 29134 3724 29178
rect 4992 29135 5044 29187
rect 3853 29047 4257 29073
rect 5034 29038 5060 29096
rect 2683 28949 2727 29007
rect 5213 29038 5239 29096
rect 14721 29038 14747 29096
rect 16236 29198 16280 29242
rect 14916 29135 14968 29187
rect 16236 29134 16280 29178
rect 14900 29038 14926 29096
rect 15703 29047 16107 29073
rect 2619 28859 2663 28917
rect 5175 28908 5815 28997
rect 14145 28908 14785 28997
rect 17233 28949 17277 29007
rect 17297 37534 17341 37592
rect 17297 28859 17341 28917
rect 17361 37198 17405 37256
rect 2555 27449 2599 27507
rect 17361 27449 17405 27507
rect 17425 37134 17469 37192
rect 2491 27359 2535 27417
rect 17425 27359 17469 27417
rect 17489 36798 17533 36856
rect 2427 25949 2471 26007
rect 17489 25949 17533 26007
rect 17553 36734 17597 36792
rect 2363 25859 2407 25917
rect 17553 25859 17597 25917
rect 17617 36597 17661 36655
rect 2299 24449 2343 24507
rect 17617 24449 17661 24507
rect 17681 36533 17725 36591
rect 2235 24359 2279 24417
rect 17681 24359 17725 24417
rect 17745 35998 17789 36056
rect 2171 22949 2215 23007
rect 17745 22949 17789 23007
rect 17809 35934 17853 35992
rect 2107 22859 2151 22917
rect 17809 22859 17853 22917
rect 17873 35598 17917 35656
rect 2043 21449 2087 21507
rect 17873 21449 17917 21507
rect 17937 35534 17981 35592
rect 1979 21359 2023 21417
rect 17937 21359 17981 21417
rect 18001 35198 18045 35256
rect 5175 21105 5815 21295
rect 14145 21105 14785 21295
rect 1915 19949 1959 20007
rect 18001 19949 18045 20007
rect 18065 35134 18109 35192
rect 1851 19859 1895 19917
rect 18065 19859 18109 19917
rect 18129 34795 18173 34853
rect 10970 19340 11090 19460
rect 10593 19066 10646 19277
rect 11002 19060 11037 19270
rect 11117 19063 11171 19273
rect 1787 18449 1831 18507
rect 18129 18449 18173 18507
rect 18193 34731 18237 34789
rect 1723 18359 1767 18417
rect 18193 18359 18237 18417
rect 18257 34398 18301 34456
rect 1659 16949 1703 17007
rect 18257 16949 18301 17007
rect 18321 34334 18365 34392
rect 1595 16859 1639 16917
rect 18321 16859 18365 16917
rect 18385 33998 18429 34056
rect 1531 15449 1575 15507
rect 18385 15449 18429 15507
rect 18449 33934 18493 33992
rect 1467 15359 1511 15417
rect 18449 15359 18493 15417
rect 18513 33598 18557 33656
rect 1403 13949 1447 14007
rect 18513 13949 18557 14007
rect 18577 33534 18621 33592
rect 1339 13859 1383 13917
rect 18577 13859 18621 13917
rect 18641 33198 18685 33256
rect 1275 12449 1319 12507
rect 18641 12449 18685 12507
rect 18705 33134 18749 33192
rect 1211 12359 1255 12417
rect 18705 12359 18749 12417
rect 18769 32798 18813 32856
rect 1147 10949 1191 11007
rect 18769 10949 18813 11007
rect 18833 32734 18877 32792
rect 1083 10859 1127 10917
rect 18833 10859 18877 10917
rect 18897 32398 18941 32456
rect 1019 9449 1063 9507
rect 18897 9449 18941 9507
rect 18961 32334 19005 32392
rect 955 9359 999 9417
rect 18961 9359 19005 9417
rect 19025 32091 19069 32149
rect 891 7949 935 8007
rect 19025 7949 19069 8007
rect 19089 32027 19133 32085
rect 827 7859 871 7917
rect 19089 7859 19133 7917
rect 19153 31598 19197 31656
rect 763 6449 807 6507
rect 19153 6449 19197 6507
rect 19217 31534 19261 31592
rect 699 6359 743 6417
rect 19217 6359 19261 6417
rect 19281 31198 19325 31256
rect 12871 6107 12965 6201
rect 12871 5483 12965 5577
rect 13009 5939 13103 6033
rect 13009 5483 13103 5577
rect 13147 5771 13241 5865
rect 13147 5483 13241 5577
rect 13285 5603 13379 5697
rect 13285 5483 13379 5577
rect 635 4949 679 5007
rect 19281 4949 19325 5007
rect 19345 31134 19389 31192
rect 571 4859 615 4917
rect 19345 4859 19389 4917
rect 19409 30798 19453 30856
rect 507 3449 551 3507
rect 19409 3449 19453 3507
rect 19473 30734 19517 30792
rect 443 3359 487 3417
rect 19473 3359 19517 3417
rect 19537 30597 19581 30655
rect 379 1949 423 2007
rect 6814 2130 6866 2156
rect 7614 2130 7666 2156
rect 8414 2130 8466 2156
rect 9214 2130 9266 2156
rect 10014 2130 10066 2156
rect 10814 2130 10866 2156
rect 11614 2130 11666 2156
rect 6086 2023 6138 2049
rect 6486 2023 6538 2049
rect 6886 2023 6938 2049
rect 7286 2023 7338 2049
rect 7686 2023 7738 2049
rect 8086 2023 8138 2049
rect 8486 2023 8538 2049
rect 8886 2023 8938 2049
rect 9286 2023 9338 2049
rect 9686 2023 9738 2049
rect 10086 2023 10138 2049
rect 10486 2023 10538 2049
rect 10886 2023 10938 2049
rect 11286 2023 11338 2049
rect 11686 2023 11738 2049
rect 12086 2023 12138 2049
rect 6814 1951 6866 1977
rect 7614 1951 7666 1977
rect 8414 1951 8466 1977
rect 9214 1951 9266 1977
rect 10014 1951 10066 1977
rect 10814 1951 10866 1977
rect 11614 1951 11666 1977
rect 315 1859 359 1917
rect 12443 1903 12517 1977
rect 19537 1949 19581 2007
rect 19601 30533 19645 30591
rect 6086 1844 6138 1870
rect 6183 1802 6235 1854
rect 6486 1844 6538 1870
rect 6583 1802 6635 1854
rect 6886 1844 6938 1870
rect 6983 1802 7035 1854
rect 7286 1844 7338 1870
rect 7383 1802 7435 1854
rect 7686 1844 7738 1870
rect 7783 1802 7835 1854
rect 8086 1844 8138 1870
rect 8183 1802 8235 1854
rect 8486 1844 8538 1870
rect 8583 1802 8635 1854
rect 8886 1844 8938 1870
rect 8983 1802 9035 1854
rect 9286 1844 9338 1870
rect 9383 1802 9435 1854
rect 9686 1844 9738 1870
rect 9783 1802 9835 1854
rect 10086 1844 10138 1870
rect 10183 1802 10235 1854
rect 10486 1844 10538 1870
rect 10583 1802 10635 1854
rect 10886 1844 10938 1870
rect 10983 1802 11035 1854
rect 11286 1844 11338 1870
rect 11383 1802 11435 1854
rect 11686 1844 11738 1870
rect 11783 1802 11835 1854
rect 12086 1844 12138 1870
rect 19601 1859 19645 1917
rect 19665 29998 19709 30056
rect 12183 1802 12235 1854
rect 6090 593 6116 987
rect 6490 593 6516 987
rect 6890 593 6916 987
rect 7290 593 7316 987
rect 7690 593 7716 987
rect 8090 593 8116 987
rect 8490 593 8516 987
rect 8890 593 8916 987
rect 9290 593 9316 987
rect 9690 593 9716 987
rect 10090 593 10116 987
rect 10490 593 10516 987
rect 10890 593 10916 987
rect 11290 593 11316 987
rect 11690 593 11716 987
rect 12090 593 12116 987
rect 251 449 295 507
rect 187 359 231 417
rect 1092 233 1136 277
rect -18215 -75 -18145 -5
rect -16215 -75 -16145 -5
rect -14215 -75 -14145 -5
rect -12215 -75 -12145 -5
rect -10215 -75 -10145 -5
rect -8215 -75 -8145 -5
rect -6215 -75 -6145 -5
rect -4215 -75 -4145 -5
rect -2215 -75 -2145 -5
rect -215 -75 -145 -5
rect -18265 -1010 -18239 -984
rect -16265 -918 -16239 -892
rect -18011 -964 -17985 -938
rect -14265 -826 -14239 -800
rect -16011 -872 -15985 -846
rect -12265 -734 -12239 -708
rect -14011 -780 -13985 -754
rect -10265 -642 -10239 -616
rect -12011 -688 -11985 -662
rect -8265 -550 -8239 -524
rect -10011 -596 -9985 -570
rect -6265 -458 -6239 -432
rect -8011 -504 -7985 -478
rect -4265 -366 -4239 -340
rect -6011 -412 -5985 -386
rect -2265 -274 -2239 -248
rect -4011 -320 -3985 -294
rect -265 -182 -239 -156
rect -2011 -228 -1985 -202
rect 1030 -90 1056 -64
rect -11 -136 15 -110
rect 7284 140 7310 166
rect 6284 48 6310 74
rect 6030 2 6056 28
rect 1284 -44 1310 -18
rect 7030 94 7056 120
rect 7450 140 7476 166
rect 7396 94 7422 120
rect 7850 48 7876 74
rect 7796 2 7822 28
rect 8250 -44 8276 -18
rect 8196 -90 8222 -64
rect 19665 449 19709 507
rect 19729 29934 19773 29992
rect 19729 359 19773 417
rect 20105 -75 20175 -5
rect 22105 -75 22175 -5
rect 24105 -75 24175 -5
rect 26105 -75 26175 -5
rect 28105 -75 28175 -5
rect 30105 -75 30175 -5
rect 32105 -75 32175 -5
rect 34105 -75 34175 -5
rect 36105 -75 36175 -5
rect 38105 -75 38175 -5
rect 12250 -136 12276 -110
rect 19944 -136 19970 -110
rect 12196 -182 12222 -156
rect 11850 -228 11876 -202
rect 11796 -274 11822 -248
rect 11450 -320 11476 -294
rect 11396 -366 11422 -340
rect 11050 -412 11076 -386
rect 10996 -458 11022 -432
rect 10650 -504 10676 -478
rect 10596 -550 10622 -524
rect 10250 -596 10276 -570
rect 10196 -642 10222 -616
rect 9850 -688 9876 -662
rect 9796 -734 9822 -708
rect 9450 -780 9476 -754
rect 9396 -826 9422 -800
rect 9050 -872 9076 -846
rect 8996 -918 9022 -892
rect 8650 -964 8676 -938
rect 8596 -1010 8622 -984
rect 20198 -182 20224 -156
rect 21944 -228 21970 -202
rect 22198 -274 22224 -248
rect 23944 -320 23970 -294
rect 24198 -366 24224 -340
rect 25944 -412 25970 -386
rect 26198 -458 26224 -432
rect 27944 -504 27970 -478
rect 28198 -550 28224 -524
rect 29944 -596 29970 -570
rect 30198 -642 30224 -616
rect 31944 -688 31970 -662
rect 32198 -734 32224 -708
rect 33944 -780 33970 -754
rect 34198 -826 34224 -800
rect 35944 -872 35970 -846
rect 36198 -918 36224 -892
rect 37944 -964 37970 -938
rect 38198 -1010 38224 -984
rect 7092 -1095 7136 -1031
rect -17940 -1220 -17820 -1100
rect -15940 -1220 -15820 -1100
rect -13940 -1220 -13820 -1100
rect -11940 -1220 -11820 -1100
rect -9940 -1220 -9820 -1100
rect -7940 -1220 -7820 -1100
rect -5940 -1220 -5820 -1100
rect -3940 -1220 -3820 -1100
rect -1940 -1220 -1820 -1100
rect 60 -1220 180 -1100
rect 1355 -1220 1475 -1100
rect 6355 -1220 6475 -1100
rect 7355 -1220 7475 -1100
rect 19776 -1220 19896 -1100
rect 21776 -1220 21896 -1100
rect 23776 -1220 23896 -1100
rect 25776 -1220 25896 -1100
rect 27776 -1220 27896 -1100
rect 29776 -1220 29896 -1100
rect 31776 -1220 31896 -1100
rect 33776 -1220 33896 -1100
rect 35776 -1220 35896 -1100
rect 37776 -1220 37896 -1100
rect -18438 -1830 -18318 -1710
rect -16438 -1830 -16318 -1710
rect -14438 -1830 -14318 -1710
rect -12438 -1830 -12318 -1710
rect -10438 -1830 -10318 -1710
rect -8438 -1830 -8318 -1710
rect -6438 -1830 -6318 -1710
rect -4438 -1830 -4318 -1710
rect -2438 -1830 -2318 -1710
rect -438 -1830 -318 -1710
rect 857 -1830 977 -1710
rect 5857 -1830 5977 -1710
rect 6857 -1830 6977 -1710
rect 20260 -1830 20380 -1710
rect 22260 -1830 22380 -1710
rect 24260 -1830 24380 -1710
rect 26260 -1830 26380 -1710
rect 28260 -1830 28380 -1710
rect 30260 -1830 30380 -1710
rect 32260 -1830 32380 -1710
rect 34260 -1830 34380 -1710
rect 36260 -1830 36380 -1710
rect 38260 -1830 38380 -1710
rect 4410 -2190 4790 -2010
rect 17220 -2180 17780 -2020
<< metal2 >>
rect 40 44259 3060 44262
rect 40 44215 2863 44259
rect 3055 44215 3060 44259
rect 40 44212 3060 44215
rect 39960 44212 40160 44262
rect 3256 44021 3306 44024
rect 3256 44010 3259 44021
rect 40 43963 3259 44010
rect 3303 43963 3306 44021
rect 40 43960 3306 43963
rect 16654 44021 16704 44024
rect 16654 43963 16657 44021
rect 16701 44010 16704 44021
rect 16701 43963 19920 44010
rect 16654 43960 19920 43963
rect 3320 43931 3370 43934
rect 3320 43920 3323 43931
rect 40 43873 3323 43920
rect 3367 43873 3370 43931
rect 40 43870 3370 43873
rect 16590 43931 16640 43934
rect 16590 43873 16593 43931
rect 16637 43920 16640 43931
rect 16637 43873 19920 43920
rect 16590 43870 19920 43873
rect 40 43817 440 43820
rect 40 43733 43 43817
rect 435 43733 440 43817
rect 40 43730 440 43733
rect 19518 43817 19920 43820
rect 19518 43733 19523 43817
rect 19915 43733 19920 43817
rect 19518 43730 19920 43733
rect 8770 42867 11190 42872
rect 8770 42777 10923 42867
rect 11113 42777 11190 42867
rect 8770 42772 11190 42777
rect 40060 42762 40160 44212
rect 40 42759 3060 42762
rect 40 42715 2863 42759
rect 3055 42715 3060 42759
rect 40 42712 3060 42715
rect 8770 42729 11190 42734
rect 8770 42639 10655 42729
rect 10845 42639 11190 42729
rect 39960 42712 40160 42762
rect 8770 42634 11190 42639
rect 8770 42591 11190 42596
rect 3384 42521 3434 42524
rect 3384 42510 3387 42521
rect 40 42463 3387 42510
rect 3431 42463 3434 42521
rect 8770 42501 10387 42591
rect 10577 42501 11190 42591
rect 8770 42496 11190 42501
rect 16526 42521 16576 42524
rect 40 42460 3434 42463
rect 16526 42463 16529 42521
rect 16573 42510 16576 42521
rect 16573 42463 19920 42510
rect 16526 42460 19920 42463
rect 8770 42453 11190 42458
rect 3448 42431 3498 42434
rect 3448 42420 3451 42431
rect 40 42373 3451 42420
rect 3495 42373 3498 42431
rect 40 42370 3498 42373
rect 8770 42363 10119 42453
rect 10309 42363 11190 42453
rect 16462 42431 16512 42434
rect 16462 42373 16465 42431
rect 16509 42420 16512 42431
rect 16509 42373 19920 42420
rect 16462 42370 19920 42373
rect 8770 42358 11190 42363
rect 40 42317 440 42320
rect 40 42233 43 42317
rect 435 42233 440 42317
rect 40 42230 440 42233
rect 8770 42315 11190 42320
rect 8770 42225 9851 42315
rect 10041 42225 11190 42315
rect 19518 42317 19920 42320
rect 19518 42233 19523 42317
rect 19915 42233 19920 42317
rect 19518 42230 19920 42233
rect 8770 42220 11190 42225
rect 5087 41793 5090 41871
rect 5170 41793 5320 41871
rect 14640 41793 14790 41871
rect 14870 41793 14873 41871
rect 3256 41642 3727 41645
rect 3256 41584 3259 41642
rect 3303 41598 3680 41642
rect 3724 41598 3727 41642
rect 3303 41595 3727 41598
rect 16233 41642 16704 41645
rect 16233 41598 16236 41642
rect 16280 41598 16657 41642
rect 16233 41595 16657 41598
rect 3303 41584 3306 41595
rect 3256 41581 3306 41584
rect 4989 41587 5190 41590
rect 3320 41578 3727 41581
rect 3320 41520 3323 41578
rect 3367 41534 3680 41578
rect 3724 41534 3727 41578
rect 3367 41531 3727 41534
rect 4989 41535 4992 41587
rect 5044 41535 5190 41587
rect 4989 41532 5190 41535
rect 14770 41587 14971 41590
rect 14770 41535 14916 41587
rect 14968 41535 14971 41587
rect 16654 41584 16657 41595
rect 16701 41584 16704 41642
rect 16654 41581 16704 41584
rect 14770 41532 14971 41535
rect 16233 41578 16640 41581
rect 16233 41534 16236 41578
rect 16280 41534 16593 41578
rect 16233 41531 16593 41534
rect 3367 41520 3370 41531
rect 3320 41517 3370 41520
rect 16590 41520 16593 41531
rect 16637 41520 16640 41578
rect 16590 41517 16640 41520
rect 5031 41496 5242 41499
rect 3850 41447 3853 41473
rect 4257 41447 4260 41473
rect 40 41259 3060 41262
rect 40 41215 2863 41259
rect 3055 41215 3060 41259
rect 40 41212 3060 41215
rect 3384 41242 3727 41245
rect 3384 41184 3387 41242
rect 3431 41198 3680 41242
rect 3724 41198 3727 41242
rect 3431 41195 3727 41198
rect 3431 41184 3434 41195
rect 3384 41181 3434 41184
rect 3448 41178 3727 41181
rect 3448 41120 3451 41178
rect 3495 41134 3680 41178
rect 3724 41134 3727 41178
rect 3495 41131 3727 41134
rect 3495 41120 3498 41131
rect 3448 41117 3498 41120
rect 3850 41073 4260 41447
rect 5031 41438 5034 41496
rect 5060 41438 5213 41496
rect 5239 41438 5242 41496
rect 5031 41435 5242 41438
rect 14718 41496 14929 41499
rect 14718 41438 14721 41496
rect 14747 41438 14900 41496
rect 14926 41438 14929 41496
rect 14718 41435 14929 41438
rect 15700 41447 15703 41473
rect 16107 41447 16110 41473
rect 4989 41187 5190 41190
rect 4989 41135 4992 41187
rect 5044 41135 5190 41187
rect 4989 41132 5190 41135
rect 14770 41187 14971 41190
rect 14770 41135 14916 41187
rect 14968 41135 14971 41187
rect 14770 41132 14971 41135
rect 3850 41047 3853 41073
rect 4257 41047 4260 41073
rect 3512 41021 3562 41024
rect 3512 41010 3515 41021
rect 40 40963 3515 41010
rect 3559 40963 3562 41021
rect 40 40960 3562 40963
rect 3576 40931 3626 40934
rect 3576 40920 3579 40931
rect 40 40873 3579 40920
rect 3623 40873 3626 40931
rect 40 40870 3626 40873
rect 3512 40842 3727 40845
rect 40 40817 440 40820
rect 40 40733 43 40817
rect 435 40733 440 40817
rect 3512 40784 3515 40842
rect 3559 40798 3680 40842
rect 3724 40798 3727 40842
rect 3559 40795 3727 40798
rect 3559 40784 3562 40795
rect 3512 40781 3562 40784
rect 40 40730 440 40733
rect 3576 40778 3727 40781
rect 3576 40720 3579 40778
rect 3623 40734 3680 40778
rect 3724 40734 3727 40778
rect 3623 40731 3727 40734
rect 3623 40720 3626 40731
rect 3576 40717 3626 40720
rect 3850 40673 4260 41047
rect 5031 41096 5242 41099
rect 5031 41038 5034 41096
rect 5060 41038 5213 41096
rect 5239 41038 5242 41096
rect 5031 41035 5242 41038
rect 14718 41096 14929 41099
rect 14718 41038 14721 41096
rect 14747 41038 14900 41096
rect 14926 41038 14929 41096
rect 14718 41035 14929 41038
rect 15700 41073 16110 41447
rect 40060 41262 40160 42712
rect 16233 41242 16576 41245
rect 16233 41198 16236 41242
rect 16280 41198 16529 41242
rect 16233 41195 16529 41198
rect 16526 41184 16529 41195
rect 16573 41184 16576 41242
rect 39960 41212 40160 41262
rect 16526 41181 16576 41184
rect 16233 41178 16512 41181
rect 16233 41134 16236 41178
rect 16280 41134 16465 41178
rect 16233 41131 16465 41134
rect 16462 41120 16465 41131
rect 16509 41120 16512 41178
rect 16462 41117 16512 41120
rect 15700 41047 15703 41073
rect 16107 41047 16110 41073
rect 5138 41018 5349 41021
rect 5138 40960 5141 41018
rect 5167 40960 5320 41018
rect 5346 40960 5349 41018
rect 5138 40957 5349 40960
rect 14611 41018 14822 41021
rect 14611 40960 14614 41018
rect 14640 40960 14793 41018
rect 14819 40960 14822 41018
rect 14611 40957 14822 40960
rect 4989 40787 5190 40790
rect 4989 40735 4992 40787
rect 5044 40735 5190 40787
rect 4989 40732 5190 40735
rect 14770 40787 14971 40790
rect 14770 40735 14916 40787
rect 14968 40735 14971 40787
rect 14770 40732 14971 40735
rect 3850 40647 3853 40673
rect 4257 40647 4260 40673
rect 3576 40456 3626 40459
rect 3576 40398 3579 40456
rect 3623 40445 3626 40456
rect 3623 40442 3727 40445
rect 3623 40398 3680 40442
rect 3724 40398 3727 40442
rect 3576 40395 3727 40398
rect 3512 40392 3562 40395
rect 3512 40334 3515 40392
rect 3559 40381 3562 40392
rect 3559 40378 3727 40381
rect 3559 40334 3680 40378
rect 3724 40334 3727 40378
rect 3512 40331 3727 40334
rect 3850 40273 4260 40647
rect 5031 40696 5242 40699
rect 5031 40638 5034 40696
rect 5060 40638 5213 40696
rect 5239 40638 5242 40696
rect 5031 40635 5242 40638
rect 14718 40696 14929 40699
rect 14718 40638 14721 40696
rect 14747 40638 14900 40696
rect 14926 40638 14929 40696
rect 14718 40635 14929 40638
rect 15700 40673 16110 41047
rect 16398 41021 16448 41024
rect 16398 40963 16401 41021
rect 16445 41010 16448 41021
rect 16445 40963 19920 41010
rect 16398 40960 19920 40963
rect 16334 40931 16384 40934
rect 16334 40873 16337 40931
rect 16381 40920 16384 40931
rect 16381 40873 19920 40920
rect 16334 40870 19920 40873
rect 16233 40842 16448 40845
rect 16233 40798 16236 40842
rect 16280 40798 16401 40842
rect 16233 40795 16401 40798
rect 16398 40784 16401 40795
rect 16445 40784 16448 40842
rect 16398 40781 16448 40784
rect 19518 40817 19920 40820
rect 16233 40778 16384 40781
rect 16233 40734 16236 40778
rect 16280 40734 16337 40778
rect 16233 40731 16337 40734
rect 16334 40720 16337 40731
rect 16381 40720 16384 40778
rect 19518 40733 19523 40817
rect 19915 40733 19920 40817
rect 19518 40730 19920 40733
rect 16334 40717 16384 40720
rect 15700 40647 15703 40673
rect 16107 40647 16110 40673
rect 4989 40387 5190 40390
rect 4989 40335 4992 40387
rect 5044 40335 5190 40387
rect 4989 40332 5190 40335
rect 14770 40387 14971 40390
rect 14770 40335 14916 40387
rect 14968 40335 14971 40387
rect 14770 40332 14971 40335
rect 3850 40247 3853 40273
rect 4257 40247 4260 40273
rect 3448 40056 3498 40059
rect 3448 39998 3451 40056
rect 3495 40045 3498 40056
rect 3495 40042 3727 40045
rect 3495 39998 3680 40042
rect 3724 39998 3727 40042
rect 3448 39995 3727 39998
rect 3384 39992 3434 39995
rect 3384 39934 3387 39992
rect 3431 39981 3434 39992
rect 3431 39978 3727 39981
rect 3431 39934 3680 39978
rect 3724 39934 3727 39978
rect 3384 39931 3727 39934
rect 3850 39873 4260 40247
rect 5031 40296 5242 40299
rect 5031 40238 5034 40296
rect 5060 40238 5213 40296
rect 5239 40238 5242 40296
rect 5031 40235 5242 40238
rect 14718 40296 14929 40299
rect 14718 40238 14721 40296
rect 14747 40238 14900 40296
rect 14926 40238 14929 40296
rect 14718 40235 14929 40238
rect 15700 40273 16110 40647
rect 16334 40456 16384 40459
rect 16334 40445 16337 40456
rect 16233 40442 16337 40445
rect 16233 40398 16236 40442
rect 16280 40398 16337 40442
rect 16381 40398 16384 40456
rect 16233 40395 16384 40398
rect 16398 40392 16448 40395
rect 16398 40381 16401 40392
rect 16233 40378 16401 40381
rect 16233 40334 16236 40378
rect 16280 40334 16401 40378
rect 16445 40334 16448 40392
rect 16233 40331 16448 40334
rect 15700 40247 15703 40273
rect 16107 40247 16110 40273
rect 5138 40218 5349 40221
rect 5138 40160 5141 40218
rect 5167 40160 5320 40218
rect 5346 40160 5349 40218
rect 5138 40157 5349 40160
rect 14611 40218 14822 40221
rect 14611 40160 14614 40218
rect 14640 40160 14793 40218
rect 14819 40160 14822 40218
rect 14611 40157 14822 40160
rect 4989 39987 5190 39990
rect 4989 39935 4992 39987
rect 5044 39935 5190 39987
rect 4989 39932 5190 39935
rect 14770 39987 14971 39990
rect 14770 39935 14916 39987
rect 14968 39935 14971 39987
rect 14770 39932 14971 39935
rect 3850 39847 3853 39873
rect 4257 39847 4260 39873
rect 40 39759 3060 39762
rect 40 39715 2863 39759
rect 3055 39715 3060 39759
rect 40 39712 3060 39715
rect 3320 39656 3370 39659
rect 3320 39598 3323 39656
rect 3367 39645 3370 39656
rect 3367 39642 3727 39645
rect 3367 39598 3680 39642
rect 3724 39598 3727 39642
rect 3320 39595 3727 39598
rect 3256 39592 3306 39595
rect 3256 39534 3259 39592
rect 3303 39581 3306 39592
rect 3303 39578 3727 39581
rect 3303 39534 3680 39578
rect 3724 39534 3727 39578
rect 3256 39531 3727 39534
rect 40 39507 3626 39510
rect 40 39460 3579 39507
rect 3576 39449 3579 39460
rect 3623 39449 3626 39507
rect 3576 39446 3626 39449
rect 3850 39473 4260 39847
rect 5031 39896 5242 39899
rect 5031 39838 5034 39896
rect 5060 39838 5213 39896
rect 5239 39838 5242 39896
rect 5031 39835 5242 39838
rect 14718 39896 14929 39899
rect 14718 39838 14721 39896
rect 14747 39838 14900 39896
rect 14926 39838 14929 39896
rect 14718 39835 14929 39838
rect 15700 39873 16110 40247
rect 16462 40056 16512 40059
rect 16462 40045 16465 40056
rect 16233 40042 16465 40045
rect 16233 39998 16236 40042
rect 16280 39998 16465 40042
rect 16509 39998 16512 40056
rect 16233 39995 16512 39998
rect 16526 39992 16576 39995
rect 16526 39981 16529 39992
rect 16233 39978 16529 39981
rect 16233 39934 16236 39978
rect 16280 39934 16529 39978
rect 16573 39934 16576 39992
rect 16233 39931 16576 39934
rect 15700 39847 15703 39873
rect 16107 39847 16110 39873
rect 4989 39587 5190 39590
rect 4989 39535 4992 39587
rect 5044 39535 5190 39587
rect 4989 39532 5190 39535
rect 14770 39587 14971 39590
rect 14770 39535 14916 39587
rect 14968 39535 14971 39587
rect 14770 39532 14971 39535
rect 3850 39447 3853 39473
rect 4257 39447 4260 39473
rect 40 39417 3562 39420
rect 40 39370 3515 39417
rect 3512 39359 3515 39370
rect 3559 39359 3562 39417
rect 3512 39356 3562 39359
rect 40 39317 440 39320
rect 40 39233 43 39317
rect 435 39233 440 39317
rect 40 39230 440 39233
rect 3192 39256 3242 39259
rect 3192 39198 3195 39256
rect 3239 39245 3242 39256
rect 3239 39242 3727 39245
rect 3239 39198 3680 39242
rect 3724 39198 3727 39242
rect 3192 39195 3727 39198
rect 3128 39192 3178 39195
rect 3128 39134 3131 39192
rect 3175 39181 3178 39192
rect 3175 39178 3727 39181
rect 3175 39134 3680 39178
rect 3724 39134 3727 39178
rect 3128 39131 3727 39134
rect 3850 39073 4260 39447
rect 5031 39496 5242 39499
rect 5031 39438 5034 39496
rect 5060 39438 5213 39496
rect 5239 39438 5242 39496
rect 5031 39435 5242 39438
rect 14718 39496 14929 39499
rect 14718 39438 14721 39496
rect 14747 39438 14900 39496
rect 14926 39438 14929 39496
rect 14718 39435 14929 39438
rect 15700 39473 16110 39847
rect 40060 39762 40160 41212
rect 39960 39712 40160 39762
rect 16590 39656 16640 39659
rect 16590 39645 16593 39656
rect 16233 39642 16593 39645
rect 16233 39598 16236 39642
rect 16280 39598 16593 39642
rect 16637 39598 16640 39656
rect 16233 39595 16640 39598
rect 16654 39592 16704 39595
rect 16654 39581 16657 39592
rect 16233 39578 16657 39581
rect 16233 39534 16236 39578
rect 16280 39534 16657 39578
rect 16701 39534 16704 39592
rect 16233 39531 16704 39534
rect 15700 39447 15703 39473
rect 16107 39447 16110 39473
rect 5138 39418 5349 39421
rect 5138 39360 5141 39418
rect 5167 39360 5320 39418
rect 5346 39360 5349 39418
rect 5138 39357 5349 39360
rect 14611 39418 14822 39421
rect 14611 39360 14614 39418
rect 14640 39360 14793 39418
rect 14819 39360 14822 39418
rect 14611 39357 14822 39360
rect 4989 39187 5190 39190
rect 4989 39135 4992 39187
rect 5044 39135 5190 39187
rect 4989 39132 5190 39135
rect 14770 39187 14971 39190
rect 14770 39135 14916 39187
rect 14968 39135 14971 39187
rect 14770 39132 14971 39135
rect 3850 39047 3853 39073
rect 4257 39047 4260 39073
rect 3064 38856 3114 38859
rect 3064 38798 3067 38856
rect 3111 38845 3114 38856
rect 3111 38842 3727 38845
rect 3111 38798 3680 38842
rect 3724 38798 3727 38842
rect 3064 38795 3727 38798
rect 3000 38792 3050 38795
rect 3000 38734 3003 38792
rect 3047 38781 3050 38792
rect 3047 38778 3727 38781
rect 3047 38734 3680 38778
rect 3724 38734 3727 38778
rect 3000 38731 3727 38734
rect 3850 38673 4260 39047
rect 5031 39096 5242 39099
rect 5031 39038 5034 39096
rect 5060 39038 5213 39096
rect 5239 39038 5242 39096
rect 5031 39035 5242 39038
rect 14718 39096 14929 39099
rect 14718 39038 14721 39096
rect 14747 39038 14900 39096
rect 14926 39038 14929 39096
rect 14718 39035 14929 39038
rect 15700 39073 16110 39447
rect 16334 39507 19920 39510
rect 16334 39449 16337 39507
rect 16381 39460 19920 39507
rect 16381 39449 16384 39460
rect 16334 39446 16384 39449
rect 16398 39417 19920 39420
rect 16398 39359 16401 39417
rect 16445 39370 19920 39417
rect 16445 39359 16448 39370
rect 16398 39356 16448 39359
rect 19518 39317 19920 39320
rect 16718 39256 16768 39259
rect 16718 39245 16721 39256
rect 16233 39242 16721 39245
rect 16233 39198 16236 39242
rect 16280 39198 16721 39242
rect 16765 39198 16768 39256
rect 19518 39233 19523 39317
rect 19915 39233 19920 39317
rect 19518 39230 19920 39233
rect 16233 39195 16768 39198
rect 16782 39192 16832 39195
rect 16782 39181 16785 39192
rect 16233 39178 16785 39181
rect 16233 39134 16236 39178
rect 16280 39134 16785 39178
rect 16829 39134 16832 39192
rect 16233 39131 16832 39134
rect 15700 39047 15703 39073
rect 16107 39047 16110 39073
rect 4989 38787 5190 38790
rect 4989 38735 4992 38787
rect 5044 38735 5190 38787
rect 4989 38732 5190 38735
rect 14770 38787 14971 38790
rect 14770 38735 14916 38787
rect 14968 38735 14971 38787
rect 14770 38732 14971 38735
rect 3850 38647 3853 38673
rect 4257 38647 4260 38673
rect 2936 38456 2986 38459
rect 2936 38398 2939 38456
rect 2983 38445 2986 38456
rect 2983 38442 3727 38445
rect 2983 38398 3680 38442
rect 3724 38398 3727 38442
rect 2936 38395 3727 38398
rect 2872 38392 2922 38395
rect 2872 38334 2875 38392
rect 2919 38381 2922 38392
rect 2919 38378 3727 38381
rect 2919 38334 3680 38378
rect 3724 38334 3727 38378
rect 2872 38331 3727 38334
rect 3850 38273 4260 38647
rect 5031 38696 5242 38699
rect 5031 38638 5034 38696
rect 5060 38638 5213 38696
rect 5239 38638 5242 38696
rect 5031 38635 5242 38638
rect 14718 38696 14929 38699
rect 14718 38638 14721 38696
rect 14747 38638 14900 38696
rect 14926 38638 14929 38696
rect 14718 38635 14929 38638
rect 15700 38673 16110 39047
rect 16846 38856 16896 38859
rect 16846 38845 16849 38856
rect 16233 38842 16849 38845
rect 16233 38798 16236 38842
rect 16280 38798 16849 38842
rect 16893 38798 16896 38856
rect 16233 38795 16896 38798
rect 16910 38792 16960 38795
rect 16910 38781 16913 38792
rect 16233 38778 16913 38781
rect 16233 38734 16236 38778
rect 16280 38734 16913 38778
rect 16957 38734 16960 38792
rect 16233 38731 16960 38734
rect 15700 38647 15703 38673
rect 16107 38647 16110 38673
rect 5138 38618 5349 38621
rect 5138 38560 5141 38618
rect 5167 38560 5320 38618
rect 5346 38560 5349 38618
rect 5138 38557 5349 38560
rect 14611 38618 14822 38621
rect 14611 38560 14614 38618
rect 14640 38560 14793 38618
rect 14819 38560 14822 38618
rect 14611 38557 14822 38560
rect 4989 38387 5190 38390
rect 4989 38335 4992 38387
rect 5044 38335 5190 38387
rect 4989 38332 5190 38335
rect 14770 38387 14971 38390
rect 14770 38335 14916 38387
rect 14968 38335 14971 38387
rect 14770 38332 14971 38335
rect 40 38259 3060 38262
rect 40 38215 2863 38259
rect 3055 38215 3060 38259
rect 40 38212 3060 38215
rect 3850 38247 3853 38273
rect 4257 38247 4260 38273
rect 2808 38155 2858 38158
rect 2808 38097 2811 38155
rect 2855 38144 2858 38155
rect 2855 38097 3638 38144
rect 2808 38094 3638 38097
rect 2744 38091 2794 38094
rect 2744 38033 2747 38091
rect 2791 38080 2794 38091
rect 2791 38033 3568 38080
rect 2744 38030 3568 38033
rect 40 38007 3498 38010
rect 40 37960 3451 38007
rect 3448 37949 3451 37960
rect 3495 37949 3498 38007
rect 3448 37946 3498 37949
rect 3518 37981 3568 38030
rect 3588 38045 3638 38094
rect 3588 38042 3727 38045
rect 3588 37998 3680 38042
rect 3724 37998 3727 38042
rect 3588 37995 3727 37998
rect 3518 37978 3727 37981
rect 3518 37934 3680 37978
rect 3724 37934 3727 37978
rect 3518 37931 3727 37934
rect 40 37917 3434 37920
rect 40 37870 3387 37917
rect 3384 37859 3387 37870
rect 3431 37859 3434 37917
rect 3384 37856 3434 37859
rect 3850 37873 4260 38247
rect 5031 38296 5242 38299
rect 5031 38238 5034 38296
rect 5060 38238 5213 38296
rect 5239 38238 5242 38296
rect 5031 38235 5242 38238
rect 14718 38296 14929 38299
rect 14718 38238 14721 38296
rect 14747 38238 14900 38296
rect 14926 38238 14929 38296
rect 14718 38235 14929 38238
rect 15700 38273 16110 38647
rect 16974 38456 17024 38459
rect 16974 38445 16977 38456
rect 16233 38442 16977 38445
rect 16233 38398 16236 38442
rect 16280 38398 16977 38442
rect 17021 38398 17024 38456
rect 16233 38395 17024 38398
rect 17038 38392 17088 38395
rect 17038 38381 17041 38392
rect 16233 38378 17041 38381
rect 16233 38334 16236 38378
rect 16280 38334 17041 38378
rect 17085 38334 17088 38392
rect 16233 38331 17088 38334
rect 15700 38247 15703 38273
rect 16107 38247 16110 38273
rect 40060 38262 40160 39712
rect 4989 37987 5190 37990
rect 4989 37935 4992 37987
rect 5044 37935 5190 37987
rect 4989 37932 5190 37935
rect 14770 37987 14971 37990
rect 14770 37935 14916 37987
rect 14968 37935 14971 37987
rect 14770 37932 14971 37935
rect 3850 37847 3853 37873
rect 4257 37847 4260 37873
rect 40 37817 440 37820
rect 40 37733 43 37817
rect 435 37733 440 37817
rect 40 37730 440 37733
rect 2680 37656 2730 37659
rect 2680 37598 2683 37656
rect 2727 37645 2730 37656
rect 2727 37642 3727 37645
rect 2727 37598 3680 37642
rect 3724 37598 3727 37642
rect 2680 37595 3727 37598
rect 2616 37592 2666 37595
rect 2616 37534 2619 37592
rect 2663 37581 2666 37592
rect 2663 37578 3727 37581
rect 2663 37534 3680 37578
rect 3724 37534 3727 37578
rect 2616 37531 3727 37534
rect 3850 37473 4260 37847
rect 5031 37896 5242 37899
rect 5031 37838 5034 37896
rect 5060 37838 5213 37896
rect 5239 37838 5242 37896
rect 5031 37835 5242 37838
rect 14718 37896 14929 37899
rect 14718 37838 14721 37896
rect 14747 37838 14900 37896
rect 14926 37838 14929 37896
rect 14718 37835 14929 37838
rect 15700 37873 16110 38247
rect 39960 38212 40160 38262
rect 17102 38155 17152 38158
rect 17102 38144 17105 38155
rect 16322 38097 17105 38144
rect 17149 38097 17152 38155
rect 16322 38094 17152 38097
rect 16322 38045 16372 38094
rect 17166 38091 17216 38094
rect 17166 38080 17169 38091
rect 16233 38042 16372 38045
rect 16233 37998 16236 38042
rect 16280 37998 16372 38042
rect 16233 37995 16372 37998
rect 16392 38033 17169 38080
rect 17213 38033 17216 38091
rect 16392 38030 17216 38033
rect 16392 37981 16442 38030
rect 16233 37978 16442 37981
rect 16233 37934 16236 37978
rect 16280 37934 16442 37978
rect 16462 38007 19920 38010
rect 16462 37949 16465 38007
rect 16509 37960 19920 38007
rect 16509 37949 16512 37960
rect 16462 37946 16512 37949
rect 16233 37931 16442 37934
rect 15700 37847 15703 37873
rect 16107 37847 16110 37873
rect 16526 37917 19920 37920
rect 16526 37859 16529 37917
rect 16573 37870 19920 37917
rect 16573 37859 16576 37870
rect 16526 37856 16576 37859
rect 5138 37818 5349 37821
rect 5138 37760 5141 37818
rect 5167 37760 5320 37818
rect 5346 37760 5349 37818
rect 5138 37757 5349 37760
rect 14611 37818 14822 37821
rect 14611 37760 14614 37818
rect 14640 37760 14793 37818
rect 14819 37760 14822 37818
rect 14611 37757 14822 37760
rect 4989 37587 5190 37590
rect 4989 37535 4992 37587
rect 5044 37535 5190 37587
rect 4989 37532 5190 37535
rect 14770 37587 14971 37590
rect 14770 37535 14916 37587
rect 14968 37535 14971 37587
rect 14770 37532 14971 37535
rect 3850 37447 3853 37473
rect 4257 37447 4260 37473
rect 2552 37256 2602 37259
rect 2552 37198 2555 37256
rect 2599 37245 2602 37256
rect 2599 37242 3727 37245
rect 2599 37198 3680 37242
rect 3724 37198 3727 37242
rect 2552 37195 3727 37198
rect 2488 37192 2538 37195
rect 2488 37134 2491 37192
rect 2535 37181 2538 37192
rect 2535 37178 3727 37181
rect 2535 37134 3680 37178
rect 3724 37134 3727 37178
rect 2488 37131 3727 37134
rect 3850 37073 4260 37447
rect 5031 37496 5242 37499
rect 5031 37438 5034 37496
rect 5060 37438 5213 37496
rect 5239 37438 5242 37496
rect 5031 37435 5242 37438
rect 14718 37496 14929 37499
rect 14718 37438 14721 37496
rect 14747 37438 14900 37496
rect 14926 37438 14929 37496
rect 14718 37435 14929 37438
rect 15700 37473 16110 37847
rect 19518 37817 19920 37820
rect 19518 37733 19523 37817
rect 19915 37733 19920 37817
rect 19518 37730 19920 37733
rect 17230 37656 17280 37659
rect 17230 37645 17233 37656
rect 16233 37642 17233 37645
rect 16233 37598 16236 37642
rect 16280 37598 17233 37642
rect 17277 37598 17280 37656
rect 16233 37595 17280 37598
rect 17294 37592 17344 37595
rect 17294 37581 17297 37592
rect 16233 37578 17297 37581
rect 16233 37534 16236 37578
rect 16280 37534 17297 37578
rect 17341 37534 17344 37592
rect 16233 37531 17344 37534
rect 15700 37447 15703 37473
rect 16107 37447 16110 37473
rect 4989 37187 5190 37190
rect 4989 37135 4992 37187
rect 5044 37135 5190 37187
rect 4989 37132 5190 37135
rect 14770 37187 14971 37190
rect 14770 37135 14916 37187
rect 14968 37135 14971 37187
rect 14770 37132 14971 37135
rect 3850 37047 3853 37073
rect 4257 37047 4260 37073
rect 2250 36959 3060 36962
rect 2250 36915 2863 36959
rect 3055 36915 3060 36959
rect 2250 36912 3060 36915
rect 2250 36762 2300 36912
rect 2424 36856 2474 36859
rect 2424 36798 2427 36856
rect 2471 36845 2474 36856
rect 2471 36842 3727 36845
rect 2471 36798 3680 36842
rect 3724 36798 3727 36842
rect 2424 36795 3727 36798
rect 40 36712 2300 36762
rect 2360 36792 2410 36795
rect 2360 36734 2363 36792
rect 2407 36781 2410 36792
rect 2407 36778 3727 36781
rect 2407 36734 3680 36778
rect 3724 36734 3727 36778
rect 2360 36731 3727 36734
rect 3850 36673 4260 37047
rect 5031 37096 5242 37099
rect 5031 37038 5034 37096
rect 5060 37038 5213 37096
rect 5239 37038 5242 37096
rect 5031 37035 5242 37038
rect 14718 37096 14929 37099
rect 14718 37038 14721 37096
rect 14747 37038 14900 37096
rect 14926 37038 14929 37096
rect 14718 37035 14929 37038
rect 15700 37073 16110 37447
rect 17358 37256 17408 37259
rect 17358 37245 17361 37256
rect 16233 37242 17361 37245
rect 16233 37198 16236 37242
rect 16280 37198 17361 37242
rect 17405 37198 17408 37256
rect 16233 37195 17408 37198
rect 17422 37192 17472 37195
rect 17422 37181 17425 37192
rect 16233 37178 17425 37181
rect 16233 37134 16236 37178
rect 16280 37134 17425 37178
rect 17469 37134 17472 37192
rect 16233 37131 17472 37134
rect 15700 37047 15703 37073
rect 16107 37047 16110 37073
rect 5138 37018 5349 37021
rect 5138 36960 5141 37018
rect 5167 36960 5320 37018
rect 5346 36960 5349 37018
rect 5138 36957 5349 36960
rect 14611 37018 14822 37021
rect 14611 36960 14614 37018
rect 14640 36960 14793 37018
rect 14819 36960 14822 37018
rect 14611 36957 14822 36960
rect 4989 36787 5190 36790
rect 4989 36735 4992 36787
rect 5044 36735 5190 36787
rect 4989 36732 5190 36735
rect 14770 36787 14971 36790
rect 14770 36735 14916 36787
rect 14968 36735 14971 36787
rect 14770 36732 14971 36735
rect 2296 36655 2346 36658
rect 2296 36597 2299 36655
rect 2343 36644 2346 36655
rect 3850 36647 3853 36673
rect 4257 36647 4260 36673
rect 2343 36597 3588 36644
rect 2296 36594 3588 36597
rect 2232 36591 2282 36594
rect 2232 36533 2235 36591
rect 2279 36580 2282 36591
rect 2279 36533 3518 36580
rect 2232 36530 3518 36533
rect 40 36507 3370 36510
rect 40 36460 3323 36507
rect 3320 36449 3323 36460
rect 3367 36449 3370 36507
rect 3320 36446 3370 36449
rect 40 36417 3306 36420
rect 40 36370 3259 36417
rect 3256 36359 3259 36370
rect 3303 36359 3306 36417
rect 3256 36356 3306 36359
rect 3468 36381 3518 36530
rect 3538 36445 3588 36594
rect 3538 36442 3727 36445
rect 3538 36398 3680 36442
rect 3724 36398 3727 36442
rect 3538 36395 3727 36398
rect 3468 36378 3727 36381
rect 3468 36334 3680 36378
rect 3724 36334 3727 36378
rect 3468 36331 3727 36334
rect 40 36317 440 36320
rect 40 36233 43 36317
rect 435 36233 440 36317
rect 40 36230 440 36233
rect 3850 36273 4260 36647
rect 5031 36696 5242 36699
rect 5031 36638 5034 36696
rect 5060 36638 5213 36696
rect 5239 36638 5242 36696
rect 5031 36635 5242 36638
rect 14718 36696 14929 36699
rect 14718 36638 14721 36696
rect 14747 36638 14900 36696
rect 14926 36638 14929 36696
rect 14718 36635 14929 36638
rect 15700 36673 16110 37047
rect 17486 36856 17536 36859
rect 17486 36845 17489 36856
rect 16233 36842 17489 36845
rect 16233 36798 16236 36842
rect 16280 36798 17489 36842
rect 17533 36798 17536 36856
rect 16233 36795 17536 36798
rect 17550 36792 17600 36795
rect 17550 36781 17553 36792
rect 16233 36778 17553 36781
rect 16233 36734 16236 36778
rect 16280 36734 17553 36778
rect 17597 36734 17600 36792
rect 40060 36762 40160 38212
rect 16233 36731 17600 36734
rect 39960 36712 40160 36762
rect 15700 36647 15703 36673
rect 16107 36647 16110 36673
rect 4989 36387 5190 36390
rect 4989 36335 4992 36387
rect 5044 36335 5190 36387
rect 4989 36332 5190 36335
rect 14770 36387 14971 36390
rect 14770 36335 14916 36387
rect 14968 36335 14971 36387
rect 14770 36332 14971 36335
rect 3850 36247 3853 36273
rect 4257 36247 4260 36273
rect 2168 36056 2218 36059
rect 2168 35998 2171 36056
rect 2215 36045 2218 36056
rect 2215 36042 3727 36045
rect 2215 35998 3680 36042
rect 3724 35998 3727 36042
rect 2168 35995 3727 35998
rect 2104 35992 2154 35995
rect 2104 35934 2107 35992
rect 2151 35981 2154 35992
rect 2151 35978 3727 35981
rect 2151 35934 3680 35978
rect 3724 35934 3727 35978
rect 2104 35931 3727 35934
rect 3850 35873 4260 36247
rect 5031 36296 5242 36299
rect 5031 36238 5034 36296
rect 5060 36238 5213 36296
rect 5239 36238 5242 36296
rect 5031 36235 5242 36238
rect 14718 36296 14929 36299
rect 14718 36238 14721 36296
rect 14747 36238 14900 36296
rect 14926 36238 14929 36296
rect 14718 36235 14929 36238
rect 15700 36273 16110 36647
rect 17614 36655 17664 36658
rect 17614 36644 17617 36655
rect 16372 36597 17617 36644
rect 17661 36597 17664 36655
rect 16372 36594 17664 36597
rect 16372 36445 16422 36594
rect 17678 36591 17728 36594
rect 17678 36580 17681 36591
rect 16233 36442 16422 36445
rect 16233 36398 16236 36442
rect 16280 36398 16422 36442
rect 16233 36395 16422 36398
rect 16442 36533 17681 36580
rect 17725 36533 17728 36591
rect 16442 36530 17728 36533
rect 16442 36381 16492 36530
rect 16590 36507 19920 36510
rect 16590 36449 16593 36507
rect 16637 36460 19920 36507
rect 16637 36449 16640 36460
rect 16590 36446 16640 36449
rect 16233 36378 16492 36381
rect 16233 36334 16236 36378
rect 16280 36334 16492 36378
rect 16654 36417 19920 36420
rect 16654 36359 16657 36417
rect 16701 36370 19920 36417
rect 16701 36359 16704 36370
rect 16654 36356 16704 36359
rect 16233 36331 16492 36334
rect 15700 36247 15703 36273
rect 16107 36247 16110 36273
rect 5138 36218 5349 36221
rect 5138 36160 5141 36218
rect 5167 36160 5320 36218
rect 5346 36160 5349 36218
rect 5138 36157 5349 36160
rect 14611 36218 14822 36221
rect 14611 36160 14614 36218
rect 14640 36160 14793 36218
rect 14819 36160 14822 36218
rect 14611 36157 14822 36160
rect 4989 35987 5190 35990
rect 4989 35935 4992 35987
rect 5044 35935 5190 35987
rect 4989 35932 5190 35935
rect 14770 35987 14971 35990
rect 14770 35935 14916 35987
rect 14968 35935 14971 35987
rect 14770 35932 14971 35935
rect 3850 35847 3853 35873
rect 4257 35847 4260 35873
rect 2040 35656 2090 35659
rect 2040 35598 2043 35656
rect 2087 35645 2090 35656
rect 2087 35642 3727 35645
rect 2087 35598 3680 35642
rect 3724 35598 3727 35642
rect 2040 35595 3727 35598
rect 1976 35592 2026 35595
rect 1976 35534 1979 35592
rect 2023 35581 2026 35592
rect 2023 35578 3727 35581
rect 2023 35534 3680 35578
rect 3724 35534 3727 35578
rect 1976 35531 3727 35534
rect 3850 35473 4260 35847
rect 5031 35896 5242 35899
rect 5031 35838 5034 35896
rect 5060 35838 5213 35896
rect 5239 35838 5242 35896
rect 5031 35835 5242 35838
rect 14718 35896 14929 35899
rect 14718 35838 14721 35896
rect 14747 35838 14900 35896
rect 14926 35838 14929 35896
rect 14718 35835 14929 35838
rect 15700 35873 16110 36247
rect 19518 36317 19920 36320
rect 19518 36233 19523 36317
rect 19915 36233 19920 36317
rect 19518 36230 19920 36233
rect 17742 36056 17792 36059
rect 17742 36045 17745 36056
rect 16233 36042 17745 36045
rect 16233 35998 16236 36042
rect 16280 35998 17745 36042
rect 17789 35998 17792 36056
rect 16233 35995 17792 35998
rect 17806 35992 17856 35995
rect 17806 35981 17809 35992
rect 16233 35978 17809 35981
rect 16233 35934 16236 35978
rect 16280 35934 17809 35978
rect 17853 35934 17856 35992
rect 16233 35931 17856 35934
rect 15700 35847 15703 35873
rect 16107 35847 16110 35873
rect 4989 35587 5190 35590
rect 4989 35535 4992 35587
rect 5044 35535 5190 35587
rect 4989 35532 5190 35535
rect 14770 35587 14971 35590
rect 14770 35535 14916 35587
rect 14968 35535 14971 35587
rect 14770 35532 14971 35535
rect 3850 35447 3853 35473
rect 4257 35447 4260 35473
rect 1690 35359 3060 35362
rect 1690 35315 2863 35359
rect 3055 35315 3060 35359
rect 1690 35312 3060 35315
rect 1690 35262 1740 35312
rect 40 35212 1740 35262
rect 1912 35256 1962 35259
rect 1912 35198 1915 35256
rect 1959 35245 1962 35256
rect 1959 35242 3727 35245
rect 1959 35198 3680 35242
rect 3724 35198 3727 35242
rect 1912 35195 3727 35198
rect 1848 35192 1898 35195
rect 1848 35134 1851 35192
rect 1895 35181 1898 35192
rect 1895 35178 3727 35181
rect 1895 35134 3680 35178
rect 3724 35134 3727 35178
rect 1848 35131 3727 35134
rect 3850 35073 4260 35447
rect 5031 35496 5242 35499
rect 5031 35438 5034 35496
rect 5060 35438 5213 35496
rect 5239 35438 5242 35496
rect 5031 35435 5242 35438
rect 14718 35496 14929 35499
rect 14718 35438 14721 35496
rect 14747 35438 14900 35496
rect 14926 35438 14929 35496
rect 14718 35435 14929 35438
rect 15700 35473 16110 35847
rect 17870 35656 17920 35659
rect 17870 35645 17873 35656
rect 16233 35642 17873 35645
rect 16233 35598 16236 35642
rect 16280 35598 17873 35642
rect 17917 35598 17920 35656
rect 16233 35595 17920 35598
rect 17934 35592 17984 35595
rect 17934 35581 17937 35592
rect 16233 35578 17937 35581
rect 16233 35534 16236 35578
rect 16280 35534 17937 35578
rect 17981 35534 17984 35592
rect 16233 35531 17984 35534
rect 15700 35447 15703 35473
rect 16107 35447 16110 35473
rect 5138 35418 5349 35421
rect 5138 35360 5141 35418
rect 5167 35360 5320 35418
rect 5346 35360 5349 35418
rect 5138 35357 5349 35360
rect 14611 35418 14822 35421
rect 14611 35360 14614 35418
rect 14640 35360 14793 35418
rect 14819 35360 14822 35418
rect 14611 35357 14822 35360
rect 4989 35187 5190 35190
rect 4989 35135 4992 35187
rect 5044 35135 5190 35187
rect 4989 35132 5190 35135
rect 14770 35187 14971 35190
rect 14770 35135 14916 35187
rect 14968 35135 14971 35187
rect 14770 35132 14971 35135
rect 3850 35047 3853 35073
rect 4257 35047 4260 35073
rect 40 35007 3242 35010
rect 40 34960 3195 35007
rect 3192 34949 3195 34960
rect 3239 34949 3242 35007
rect 3192 34946 3242 34949
rect 40 34917 3178 34920
rect 40 34870 3131 34917
rect 3128 34859 3131 34870
rect 3175 34859 3178 34917
rect 3128 34856 3178 34859
rect 1784 34853 1834 34856
rect 40 34817 440 34820
rect 40 34733 43 34817
rect 435 34733 440 34817
rect 1784 34795 1787 34853
rect 1831 34842 1834 34853
rect 3193 34842 3727 34845
rect 1831 34798 3680 34842
rect 3724 34798 3727 34842
rect 1831 34795 3727 34798
rect 1784 34792 3207 34795
rect 40 34730 440 34733
rect 1720 34789 1770 34792
rect 1720 34731 1723 34789
rect 1767 34778 1770 34789
rect 3216 34778 3727 34781
rect 1767 34734 3680 34778
rect 3724 34734 3727 34778
rect 1767 34731 3727 34734
rect 1720 34728 3230 34731
rect 3850 34673 4260 35047
rect 5031 35096 5242 35099
rect 5031 35038 5034 35096
rect 5060 35038 5213 35096
rect 5239 35038 5242 35096
rect 5031 35035 5242 35038
rect 14718 35096 14929 35099
rect 14718 35038 14721 35096
rect 14747 35038 14900 35096
rect 14926 35038 14929 35096
rect 14718 35035 14929 35038
rect 15700 35073 16110 35447
rect 40060 35262 40160 36712
rect 17998 35256 18048 35259
rect 17998 35245 18001 35256
rect 16233 35242 18001 35245
rect 16233 35198 16236 35242
rect 16280 35198 18001 35242
rect 18045 35198 18048 35256
rect 39960 35212 40160 35262
rect 16233 35195 18048 35198
rect 18062 35192 18112 35195
rect 18062 35181 18065 35192
rect 16233 35178 18065 35181
rect 16233 35134 16236 35178
rect 16280 35134 18065 35178
rect 18109 35134 18112 35192
rect 16233 35131 18112 35134
rect 15700 35047 15703 35073
rect 16107 35047 16110 35073
rect 4989 34787 5190 34790
rect 4989 34735 4992 34787
rect 5044 34735 5190 34787
rect 4989 34732 5190 34735
rect 14770 34787 14971 34790
rect 14770 34735 14916 34787
rect 14968 34735 14971 34787
rect 14770 34732 14971 34735
rect 3850 34647 3853 34673
rect 4257 34647 4260 34673
rect 1656 34456 1706 34459
rect 1656 34398 1659 34456
rect 1703 34445 1706 34456
rect 1703 34442 3727 34445
rect 1703 34398 3680 34442
rect 3724 34398 3727 34442
rect 1656 34395 3727 34398
rect 1592 34392 1642 34395
rect 1592 34334 1595 34392
rect 1639 34381 1642 34392
rect 1639 34378 3727 34381
rect 1639 34334 3680 34378
rect 3724 34334 3727 34378
rect 1592 34331 3727 34334
rect 3850 34273 4260 34647
rect 5031 34696 5242 34699
rect 5031 34638 5034 34696
rect 5060 34638 5213 34696
rect 5239 34638 5242 34696
rect 5031 34635 5242 34638
rect 14718 34696 14929 34699
rect 14718 34638 14721 34696
rect 14747 34638 14900 34696
rect 14926 34638 14929 34696
rect 14718 34635 14929 34638
rect 15700 34673 16110 35047
rect 16718 35007 19920 35010
rect 16718 34949 16721 35007
rect 16765 34960 19920 35007
rect 16765 34949 16768 34960
rect 16718 34946 16768 34949
rect 16782 34917 19920 34920
rect 16782 34859 16785 34917
rect 16829 34870 19920 34917
rect 16829 34859 16832 34870
rect 16782 34856 16832 34859
rect 18126 34853 18176 34856
rect 16233 34842 16767 34845
rect 18126 34842 18129 34853
rect 16233 34798 16236 34842
rect 16280 34798 18129 34842
rect 16233 34795 18129 34798
rect 18173 34795 18176 34853
rect 16753 34792 18176 34795
rect 19518 34817 19920 34820
rect 18190 34789 18240 34792
rect 16233 34778 16744 34781
rect 18190 34778 18193 34789
rect 16233 34734 16236 34778
rect 16280 34734 18193 34778
rect 16233 34731 18193 34734
rect 18237 34731 18240 34789
rect 16730 34728 18240 34731
rect 19518 34733 19523 34817
rect 19915 34733 19920 34817
rect 19518 34730 19920 34733
rect 15700 34647 15703 34673
rect 16107 34647 16110 34673
rect 5138 34618 5349 34621
rect 5138 34560 5141 34618
rect 5167 34560 5320 34618
rect 5346 34560 5349 34618
rect 5138 34557 5349 34560
rect 14611 34618 14822 34621
rect 14611 34560 14614 34618
rect 14640 34560 14793 34618
rect 14819 34560 14822 34618
rect 14611 34557 14822 34560
rect 4989 34387 5190 34390
rect 4989 34335 4992 34387
rect 5044 34335 5190 34387
rect 4989 34332 5190 34335
rect 14770 34387 14971 34390
rect 14770 34335 14916 34387
rect 14968 34335 14971 34387
rect 14770 34332 14971 34335
rect 3850 34247 3853 34273
rect 4257 34247 4260 34273
rect 1528 34056 1578 34059
rect 1528 33998 1531 34056
rect 1575 34045 1578 34056
rect 1575 34042 3727 34045
rect 1575 33998 3680 34042
rect 3724 33998 3727 34042
rect 1528 33995 3727 33998
rect 1464 33992 1514 33995
rect 1464 33934 1467 33992
rect 1511 33981 1514 33992
rect 1511 33978 3727 33981
rect 1511 33934 3680 33978
rect 3724 33934 3727 33978
rect 1464 33931 3727 33934
rect 3850 33873 4260 34247
rect 5031 34296 5242 34299
rect 5031 34238 5034 34296
rect 5060 34238 5213 34296
rect 5239 34238 5242 34296
rect 5031 34235 5242 34238
rect 14718 34296 14929 34299
rect 14718 34238 14721 34296
rect 14747 34238 14900 34296
rect 14926 34238 14929 34296
rect 14718 34235 14929 34238
rect 15700 34273 16110 34647
rect 18254 34456 18304 34459
rect 18254 34445 18257 34456
rect 16233 34442 18257 34445
rect 16233 34398 16236 34442
rect 16280 34398 18257 34442
rect 18301 34398 18304 34456
rect 16233 34395 18304 34398
rect 18318 34392 18368 34395
rect 18318 34381 18321 34392
rect 16233 34378 18321 34381
rect 16233 34334 16236 34378
rect 16280 34334 18321 34378
rect 18365 34334 18368 34392
rect 16233 34331 18368 34334
rect 15700 34247 15703 34273
rect 16107 34247 16110 34273
rect 4989 33987 5190 33990
rect 4989 33935 4992 33987
rect 5044 33935 5190 33987
rect 4989 33932 5190 33935
rect 14770 33987 14971 33990
rect 14770 33935 14916 33987
rect 14968 33935 14971 33987
rect 14770 33932 14971 33935
rect 3850 33847 3853 33873
rect 4257 33847 4260 33873
rect 40 33759 3060 33762
rect 40 33715 2863 33759
rect 3055 33715 3060 33759
rect 40 33712 3060 33715
rect 1400 33656 1450 33659
rect 1400 33598 1403 33656
rect 1447 33645 1450 33656
rect 1447 33642 3727 33645
rect 1447 33598 3680 33642
rect 3724 33598 3727 33642
rect 1400 33595 3727 33598
rect 1336 33592 1386 33595
rect 1336 33534 1339 33592
rect 1383 33581 1386 33592
rect 1383 33578 3727 33581
rect 1383 33534 3680 33578
rect 3724 33534 3727 33578
rect 1336 33531 3727 33534
rect 40 33507 3114 33510
rect 40 33460 3067 33507
rect 3064 33449 3067 33460
rect 3111 33449 3114 33507
rect 3064 33446 3114 33449
rect 3850 33473 4260 33847
rect 5031 33896 5242 33899
rect 5031 33838 5034 33896
rect 5060 33838 5213 33896
rect 5239 33838 5242 33896
rect 5031 33835 5242 33838
rect 14718 33896 14929 33899
rect 14718 33838 14721 33896
rect 14747 33838 14900 33896
rect 14926 33838 14929 33896
rect 14718 33835 14929 33838
rect 15700 33873 16110 34247
rect 18382 34056 18432 34059
rect 18382 34045 18385 34056
rect 16233 34042 18385 34045
rect 16233 33998 16236 34042
rect 16280 33998 18385 34042
rect 18429 33998 18432 34056
rect 16233 33995 18432 33998
rect 18446 33992 18496 33995
rect 18446 33981 18449 33992
rect 16233 33978 18449 33981
rect 16233 33934 16236 33978
rect 16280 33934 18449 33978
rect 18493 33934 18496 33992
rect 16233 33931 18496 33934
rect 15700 33847 15703 33873
rect 16107 33847 16110 33873
rect 5138 33818 5349 33821
rect 5138 33760 5141 33818
rect 5167 33760 5320 33818
rect 5346 33760 5349 33818
rect 5138 33757 5349 33760
rect 14611 33818 14822 33821
rect 14611 33760 14614 33818
rect 14640 33760 14793 33818
rect 14819 33760 14822 33818
rect 14611 33757 14822 33760
rect 4989 33587 5190 33590
rect 4989 33535 4992 33587
rect 5044 33535 5190 33587
rect 4989 33532 5190 33535
rect 14770 33587 14971 33590
rect 14770 33535 14916 33587
rect 14968 33535 14971 33587
rect 14770 33532 14971 33535
rect 3850 33447 3853 33473
rect 4257 33447 4260 33473
rect 40 33417 3050 33420
rect 40 33370 3003 33417
rect 3000 33359 3003 33370
rect 3047 33359 3050 33417
rect 3000 33356 3050 33359
rect 40 33317 440 33320
rect 40 33233 43 33317
rect 435 33233 440 33317
rect 40 33230 440 33233
rect 1272 33256 1322 33259
rect 1272 33198 1275 33256
rect 1319 33245 1322 33256
rect 1319 33242 3727 33245
rect 1319 33198 3680 33242
rect 3724 33198 3727 33242
rect 1272 33195 3727 33198
rect 1208 33192 1258 33195
rect 1208 33134 1211 33192
rect 1255 33181 1258 33192
rect 1255 33178 3727 33181
rect 1255 33134 3680 33178
rect 3724 33134 3727 33178
rect 1208 33131 3727 33134
rect 3850 33073 4260 33447
rect 5031 33496 5242 33499
rect 5031 33438 5034 33496
rect 5060 33438 5213 33496
rect 5239 33438 5242 33496
rect 5031 33435 5242 33438
rect 14718 33496 14929 33499
rect 14718 33438 14721 33496
rect 14747 33438 14900 33496
rect 14926 33438 14929 33496
rect 14718 33435 14929 33438
rect 15700 33473 16110 33847
rect 40060 33762 40160 35212
rect 39960 33712 40160 33762
rect 18510 33656 18560 33659
rect 18510 33645 18513 33656
rect 16233 33642 18513 33645
rect 16233 33598 16236 33642
rect 16280 33598 18513 33642
rect 18557 33598 18560 33656
rect 16233 33595 18560 33598
rect 18574 33592 18624 33595
rect 18574 33581 18577 33592
rect 16233 33578 18577 33581
rect 16233 33534 16236 33578
rect 16280 33534 18577 33578
rect 18621 33534 18624 33592
rect 16233 33531 18624 33534
rect 15700 33447 15703 33473
rect 16107 33447 16110 33473
rect 4989 33187 5190 33190
rect 4989 33135 4992 33187
rect 5044 33135 5190 33187
rect 4989 33132 5190 33135
rect 14770 33187 14971 33190
rect 14770 33135 14916 33187
rect 14968 33135 14971 33187
rect 14770 33132 14971 33135
rect 3850 33047 3853 33073
rect 4257 33047 4260 33073
rect 1144 32856 1194 32859
rect 1144 32798 1147 32856
rect 1191 32845 1194 32856
rect 1191 32842 3727 32845
rect 1191 32798 3680 32842
rect 3724 32798 3727 32842
rect 1144 32795 3727 32798
rect 1080 32792 1130 32795
rect 1080 32734 1083 32792
rect 1127 32781 1130 32792
rect 1127 32778 3727 32781
rect 1127 32734 3680 32778
rect 3724 32734 3727 32778
rect 1080 32731 3727 32734
rect 3850 32673 4260 33047
rect 5031 33096 5242 33099
rect 5031 33038 5034 33096
rect 5060 33038 5213 33096
rect 5239 33038 5242 33096
rect 5031 33035 5242 33038
rect 14718 33096 14929 33099
rect 14718 33038 14721 33096
rect 14747 33038 14900 33096
rect 14926 33038 14929 33096
rect 14718 33035 14929 33038
rect 15700 33073 16110 33447
rect 16846 33507 19920 33510
rect 16846 33449 16849 33507
rect 16893 33460 19920 33507
rect 16893 33449 16896 33460
rect 16846 33446 16896 33449
rect 16910 33417 19920 33420
rect 16910 33359 16913 33417
rect 16957 33370 19920 33417
rect 16957 33359 16960 33370
rect 16910 33356 16960 33359
rect 19518 33317 19920 33320
rect 18638 33256 18688 33259
rect 18638 33245 18641 33256
rect 16233 33242 18641 33245
rect 16233 33198 16236 33242
rect 16280 33198 18641 33242
rect 18685 33198 18688 33256
rect 19518 33233 19523 33317
rect 19915 33233 19920 33317
rect 19518 33230 19920 33233
rect 16233 33195 18688 33198
rect 18702 33192 18752 33195
rect 18702 33181 18705 33192
rect 16233 33178 18705 33181
rect 16233 33134 16236 33178
rect 16280 33134 18705 33178
rect 18749 33134 18752 33192
rect 16233 33131 18752 33134
rect 15700 33047 15703 33073
rect 16107 33047 16110 33073
rect 5138 33018 5349 33021
rect 5138 32960 5141 33018
rect 5167 32960 5320 33018
rect 5346 32960 5349 33018
rect 5138 32957 5349 32960
rect 14611 33018 14822 33021
rect 14611 32960 14614 33018
rect 14640 32960 14793 33018
rect 14819 32960 14822 33018
rect 14611 32957 14822 32960
rect 4989 32787 5190 32790
rect 4989 32735 4992 32787
rect 5044 32735 5190 32787
rect 4989 32732 5190 32735
rect 14770 32787 14971 32790
rect 14770 32735 14916 32787
rect 14968 32735 14971 32787
rect 14770 32732 14971 32735
rect 3850 32647 3853 32673
rect 4257 32647 4260 32673
rect 1016 32456 1066 32459
rect 1016 32398 1019 32456
rect 1063 32445 1066 32456
rect 1063 32442 3727 32445
rect 1063 32398 3680 32442
rect 3724 32398 3727 32442
rect 1016 32395 3727 32398
rect 952 32392 1002 32395
rect 952 32334 955 32392
rect 999 32381 1002 32392
rect 999 32378 3727 32381
rect 999 32334 3680 32378
rect 3724 32334 3727 32378
rect 952 32331 3727 32334
rect 3850 32273 4260 32647
rect 5031 32696 5242 32699
rect 5031 32638 5034 32696
rect 5060 32638 5213 32696
rect 5239 32638 5242 32696
rect 5031 32635 5242 32638
rect 14718 32696 14929 32699
rect 14718 32638 14721 32696
rect 14747 32638 14900 32696
rect 14926 32638 14929 32696
rect 14718 32635 14929 32638
rect 15700 32673 16110 33047
rect 18766 32856 18816 32859
rect 18766 32845 18769 32856
rect 16233 32842 18769 32845
rect 16233 32798 16236 32842
rect 16280 32798 18769 32842
rect 18813 32798 18816 32856
rect 16233 32795 18816 32798
rect 18830 32792 18880 32795
rect 18830 32781 18833 32792
rect 16233 32778 18833 32781
rect 16233 32734 16236 32778
rect 16280 32734 18833 32778
rect 18877 32734 18880 32792
rect 16233 32731 18880 32734
rect 15700 32647 15703 32673
rect 16107 32647 16110 32673
rect 4989 32387 5190 32390
rect 4989 32335 4992 32387
rect 5044 32335 5190 32387
rect 4989 32332 5190 32335
rect 14770 32387 14971 32390
rect 14770 32335 14916 32387
rect 14968 32335 14971 32387
rect 14770 32332 14971 32335
rect 40 32259 3060 32262
rect 40 32215 2863 32259
rect 3055 32215 3060 32259
rect 40 32212 3060 32215
rect 3850 32247 3853 32273
rect 4257 32247 4260 32273
rect 888 32149 938 32152
rect 888 32091 891 32149
rect 935 32138 938 32149
rect 935 32091 3588 32138
rect 888 32088 3588 32091
rect 824 32085 874 32088
rect 824 32027 827 32085
rect 871 32074 874 32085
rect 871 32027 3518 32074
rect 824 32024 3518 32027
rect 40 32007 2986 32010
rect 40 31960 2939 32007
rect 2936 31949 2939 31960
rect 2983 31949 2986 32007
rect 2936 31946 2986 31949
rect 3468 31981 3518 32024
rect 3538 32045 3588 32088
rect 3538 32042 3727 32045
rect 3538 31998 3680 32042
rect 3724 31998 3727 32042
rect 3538 31995 3727 31998
rect 3468 31978 3727 31981
rect 3468 31934 3680 31978
rect 3724 31934 3727 31978
rect 3468 31931 3727 31934
rect 40 31917 2922 31920
rect 40 31870 2875 31917
rect 2872 31859 2875 31870
rect 2919 31859 2922 31917
rect 2872 31856 2922 31859
rect 3850 31873 4260 32247
rect 5031 32296 5242 32299
rect 5031 32238 5034 32296
rect 5060 32238 5213 32296
rect 5239 32238 5242 32296
rect 5031 32235 5242 32238
rect 14718 32296 14929 32299
rect 14718 32238 14721 32296
rect 14747 32238 14900 32296
rect 14926 32238 14929 32296
rect 14718 32235 14929 32238
rect 15700 32273 16110 32647
rect 18894 32456 18944 32459
rect 18894 32445 18897 32456
rect 16233 32442 18897 32445
rect 16233 32398 16236 32442
rect 16280 32398 18897 32442
rect 18941 32398 18944 32456
rect 16233 32395 18944 32398
rect 18958 32392 19008 32395
rect 18958 32381 18961 32392
rect 16233 32378 18961 32381
rect 16233 32334 16236 32378
rect 16280 32334 18961 32378
rect 19005 32334 19008 32392
rect 16233 32331 19008 32334
rect 15700 32247 15703 32273
rect 16107 32247 16110 32273
rect 40060 32262 40160 33712
rect 5138 32218 5349 32221
rect 5138 32160 5141 32218
rect 5167 32160 5320 32218
rect 5346 32160 5349 32218
rect 5138 32157 5349 32160
rect 14611 32218 14822 32221
rect 14611 32160 14614 32218
rect 14640 32160 14793 32218
rect 14819 32160 14822 32218
rect 14611 32157 14822 32160
rect 4989 31987 5190 31990
rect 4989 31935 4992 31987
rect 5044 31935 5190 31987
rect 4989 31932 5190 31935
rect 14770 31987 14971 31990
rect 14770 31935 14916 31987
rect 14968 31935 14971 31987
rect 14770 31932 14971 31935
rect 3850 31847 3853 31873
rect 4257 31847 4260 31873
rect 40 31817 440 31820
rect 40 31733 43 31817
rect 435 31733 440 31817
rect 40 31730 440 31733
rect 760 31656 810 31659
rect 760 31598 763 31656
rect 807 31645 810 31656
rect 807 31642 3727 31645
rect 807 31598 3680 31642
rect 3724 31598 3727 31642
rect 760 31595 3727 31598
rect 696 31592 746 31595
rect 696 31534 699 31592
rect 743 31581 746 31592
rect 743 31578 3727 31581
rect 743 31534 3680 31578
rect 3724 31534 3727 31578
rect 696 31531 3727 31534
rect 3850 31473 4260 31847
rect 5031 31896 5242 31899
rect 5031 31838 5034 31896
rect 5060 31838 5213 31896
rect 5239 31838 5242 31896
rect 5031 31835 5242 31838
rect 14718 31896 14929 31899
rect 14718 31838 14721 31896
rect 14747 31838 14900 31896
rect 14926 31838 14929 31896
rect 14718 31835 14929 31838
rect 15700 31873 16110 32247
rect 39960 32212 40160 32262
rect 19022 32149 19072 32152
rect 19022 32138 19025 32149
rect 16372 32091 19025 32138
rect 19069 32091 19072 32149
rect 16372 32088 19072 32091
rect 16372 32045 16422 32088
rect 19086 32085 19136 32088
rect 19086 32074 19089 32085
rect 16233 32042 16422 32045
rect 16233 31998 16236 32042
rect 16280 31998 16422 32042
rect 16233 31995 16422 31998
rect 16442 32027 19089 32074
rect 19133 32027 19136 32085
rect 16442 32024 19136 32027
rect 16442 31981 16492 32024
rect 16233 31978 16492 31981
rect 16233 31934 16236 31978
rect 16280 31934 16492 31978
rect 16974 32007 19920 32010
rect 16974 31949 16977 32007
rect 17021 31960 19920 32007
rect 17021 31949 17024 31960
rect 16974 31946 17024 31949
rect 16233 31931 16492 31934
rect 15700 31847 15703 31873
rect 16107 31847 16110 31873
rect 17038 31917 19920 31920
rect 17038 31859 17041 31917
rect 17085 31870 19920 31917
rect 17085 31859 17088 31870
rect 17038 31856 17088 31859
rect 4989 31587 5190 31590
rect 4989 31535 4992 31587
rect 5044 31535 5190 31587
rect 4989 31532 5190 31535
rect 14770 31587 14971 31590
rect 14770 31535 14916 31587
rect 14968 31535 14971 31587
rect 14770 31532 14971 31535
rect 3850 31447 3853 31473
rect 4257 31447 4260 31473
rect 632 31256 682 31259
rect 632 31198 635 31256
rect 679 31245 682 31256
rect 679 31242 3727 31245
rect 679 31198 3680 31242
rect 3724 31198 3727 31242
rect 632 31195 3727 31198
rect 568 31192 618 31195
rect 568 31134 571 31192
rect 615 31181 618 31192
rect 615 31178 3727 31181
rect 615 31134 3680 31178
rect 3724 31134 3727 31178
rect 568 31131 3727 31134
rect 3850 31073 4260 31447
rect 5031 31496 5242 31499
rect 5031 31438 5034 31496
rect 5060 31438 5213 31496
rect 5239 31438 5242 31496
rect 5031 31435 5242 31438
rect 14718 31496 14929 31499
rect 14718 31438 14721 31496
rect 14747 31438 14900 31496
rect 14926 31438 14929 31496
rect 14718 31435 14929 31438
rect 15700 31473 16110 31847
rect 19518 31817 19920 31820
rect 19518 31733 19523 31817
rect 19915 31733 19920 31817
rect 19518 31730 19920 31733
rect 19150 31656 19200 31659
rect 19150 31645 19153 31656
rect 16233 31642 19153 31645
rect 16233 31598 16236 31642
rect 16280 31598 19153 31642
rect 19197 31598 19200 31656
rect 16233 31595 19200 31598
rect 19214 31592 19264 31595
rect 19214 31581 19217 31592
rect 16233 31578 19217 31581
rect 16233 31534 16236 31578
rect 16280 31534 19217 31578
rect 19261 31534 19264 31592
rect 16233 31531 19264 31534
rect 15700 31447 15703 31473
rect 16107 31447 16110 31473
rect 5138 31418 5349 31421
rect 5138 31360 5141 31418
rect 5167 31360 5320 31418
rect 5346 31360 5349 31418
rect 5138 31357 5349 31360
rect 14611 31418 14822 31421
rect 14611 31360 14614 31418
rect 14640 31360 14793 31418
rect 14819 31360 14822 31418
rect 14611 31357 14822 31360
rect 4989 31187 5190 31190
rect 4989 31135 4992 31187
rect 5044 31135 5190 31187
rect 4989 31132 5190 31135
rect 14770 31187 14971 31190
rect 14770 31135 14916 31187
rect 14968 31135 14971 31187
rect 14770 31132 14971 31135
rect 3850 31047 3853 31073
rect 4257 31047 4260 31073
rect 350 30959 3060 30962
rect 350 30915 2863 30959
rect 3055 30915 3060 30959
rect 350 30912 3060 30915
rect 350 30762 400 30912
rect 504 30856 554 30859
rect 504 30798 507 30856
rect 551 30845 554 30856
rect 551 30842 3727 30845
rect 551 30798 3680 30842
rect 3724 30798 3727 30842
rect 504 30795 3727 30798
rect 40 30712 400 30762
rect 440 30792 490 30795
rect 440 30734 443 30792
rect 487 30781 490 30792
rect 487 30778 3727 30781
rect 487 30734 3680 30778
rect 3724 30734 3727 30778
rect 440 30731 3727 30734
rect 3850 30673 4260 31047
rect 5031 31096 5242 31099
rect 5031 31038 5034 31096
rect 5060 31038 5213 31096
rect 5239 31038 5242 31096
rect 5031 31035 5242 31038
rect 14718 31096 14929 31099
rect 14718 31038 14721 31096
rect 14747 31038 14900 31096
rect 14926 31038 14929 31096
rect 14718 31035 14929 31038
rect 15700 31073 16110 31447
rect 19278 31256 19328 31259
rect 19278 31245 19281 31256
rect 16233 31242 19281 31245
rect 16233 31198 16236 31242
rect 16280 31198 19281 31242
rect 19325 31198 19328 31256
rect 16233 31195 19328 31198
rect 19342 31192 19392 31195
rect 19342 31181 19345 31192
rect 16233 31178 19345 31181
rect 16233 31134 16236 31178
rect 16280 31134 19345 31178
rect 19389 31134 19392 31192
rect 16233 31131 19392 31134
rect 15700 31047 15703 31073
rect 16107 31047 16110 31073
rect 4989 30787 5190 30790
rect 4989 30735 4992 30787
rect 5044 30735 5190 30787
rect 4989 30732 5190 30735
rect 14770 30787 14971 30790
rect 14770 30735 14916 30787
rect 14968 30735 14971 30787
rect 14770 30732 14971 30735
rect 376 30655 426 30658
rect 376 30597 379 30655
rect 423 30644 426 30655
rect 3850 30647 3853 30673
rect 4257 30647 4260 30673
rect 423 30597 3588 30644
rect 376 30594 3588 30597
rect 312 30591 362 30594
rect 312 30533 315 30591
rect 359 30580 362 30591
rect 359 30533 3518 30580
rect 312 30530 3518 30533
rect 40 30507 2858 30510
rect 40 30460 2811 30507
rect 2808 30449 2811 30460
rect 2855 30449 2858 30507
rect 2808 30446 2858 30449
rect 40 30417 2794 30420
rect 40 30370 2747 30417
rect 2744 30359 2747 30370
rect 2791 30359 2794 30417
rect 2744 30356 2794 30359
rect 3468 30381 3518 30530
rect 3538 30445 3588 30594
rect 3538 30442 3727 30445
rect 3538 30398 3680 30442
rect 3724 30398 3727 30442
rect 3538 30395 3727 30398
rect 3468 30378 3727 30381
rect 3468 30334 3680 30378
rect 3724 30334 3727 30378
rect 3468 30331 3727 30334
rect 40 30317 440 30320
rect 40 30233 43 30317
rect 435 30233 440 30317
rect 40 30230 440 30233
rect 3850 30273 4260 30647
rect 5031 30696 5242 30699
rect 5031 30638 5034 30696
rect 5060 30638 5213 30696
rect 5239 30638 5242 30696
rect 5031 30635 5242 30638
rect 14718 30696 14929 30699
rect 14718 30638 14721 30696
rect 14747 30638 14900 30696
rect 14926 30638 14929 30696
rect 14718 30635 14929 30638
rect 15700 30673 16110 31047
rect 19406 30856 19456 30859
rect 19406 30845 19409 30856
rect 16233 30842 19409 30845
rect 16233 30798 16236 30842
rect 16280 30798 19409 30842
rect 19453 30798 19456 30856
rect 16233 30795 19456 30798
rect 19470 30792 19520 30795
rect 19470 30781 19473 30792
rect 16233 30778 19473 30781
rect 16233 30734 16236 30778
rect 16280 30734 19473 30778
rect 19517 30734 19520 30792
rect 40060 30762 40160 32212
rect 16233 30731 19520 30734
rect 39960 30712 40160 30762
rect 15700 30647 15703 30673
rect 16107 30647 16110 30673
rect 5138 30618 5349 30621
rect 5138 30560 5141 30618
rect 5167 30560 5320 30618
rect 5346 30560 5349 30618
rect 5138 30557 5349 30560
rect 14611 30618 14822 30621
rect 14611 30560 14614 30618
rect 14640 30560 14793 30618
rect 14819 30560 14822 30618
rect 14611 30557 14822 30560
rect 4989 30387 5190 30390
rect 4989 30335 4992 30387
rect 5044 30335 5190 30387
rect 4989 30332 5190 30335
rect 14770 30387 14971 30390
rect 14770 30335 14916 30387
rect 14968 30335 14971 30387
rect 14770 30332 14971 30335
rect 3850 30247 3853 30273
rect 4257 30247 4260 30273
rect 248 30056 298 30059
rect 248 29998 251 30056
rect 295 30045 298 30056
rect 295 30042 3727 30045
rect 295 29998 3680 30042
rect 3724 29998 3727 30042
rect 248 29995 3727 29998
rect 184 29992 234 29995
rect 184 29934 187 29992
rect 231 29981 234 29992
rect 231 29978 3727 29981
rect 231 29934 3680 29978
rect 3724 29934 3727 29978
rect 184 29931 3727 29934
rect 3850 29873 4260 30247
rect 5031 30296 5242 30299
rect 5031 30238 5034 30296
rect 5060 30238 5213 30296
rect 5239 30238 5242 30296
rect 5031 30235 5242 30238
rect 14718 30296 14929 30299
rect 14718 30238 14721 30296
rect 14747 30238 14900 30296
rect 14926 30238 14929 30296
rect 14718 30235 14929 30238
rect 15700 30273 16110 30647
rect 19534 30655 19584 30658
rect 19534 30644 19537 30655
rect 16372 30597 19537 30644
rect 19581 30597 19584 30655
rect 16372 30594 19584 30597
rect 16372 30445 16422 30594
rect 19598 30591 19648 30594
rect 19598 30580 19601 30591
rect 16233 30442 16422 30445
rect 16233 30398 16236 30442
rect 16280 30398 16422 30442
rect 16233 30395 16422 30398
rect 16442 30533 19601 30580
rect 19645 30533 19648 30591
rect 16442 30530 19648 30533
rect 16442 30381 16492 30530
rect 17102 30507 19920 30510
rect 17102 30449 17105 30507
rect 17149 30460 19920 30507
rect 17149 30449 17152 30460
rect 17102 30446 17152 30449
rect 16233 30378 16492 30381
rect 16233 30334 16236 30378
rect 16280 30334 16492 30378
rect 17166 30417 19920 30420
rect 17166 30359 17169 30417
rect 17213 30370 19920 30417
rect 17213 30359 17216 30370
rect 17166 30356 17216 30359
rect 16233 30331 16492 30334
rect 15700 30247 15703 30273
rect 16107 30247 16110 30273
rect 4989 29987 5190 29990
rect 4989 29935 4992 29987
rect 5044 29935 5190 29987
rect 4989 29932 5190 29935
rect 14770 29987 14971 29990
rect 14770 29935 14916 29987
rect 14968 29935 14971 29987
rect 14770 29932 14971 29935
rect 3850 29847 3853 29873
rect 4257 29847 4260 29873
rect 3677 29642 3727 29645
rect 3677 29598 3680 29642
rect 3724 29598 3727 29642
rect 3677 29595 3727 29598
rect 3677 29578 3727 29581
rect 3677 29534 3680 29578
rect 3724 29534 3727 29578
rect 3677 29531 3727 29534
rect 3850 29473 4260 29847
rect 5031 29896 5242 29899
rect 5031 29838 5034 29896
rect 5060 29838 5213 29896
rect 5239 29838 5242 29896
rect 5031 29835 5242 29838
rect 14718 29896 14929 29899
rect 14718 29838 14721 29896
rect 14747 29838 14900 29896
rect 14926 29838 14929 29896
rect 14718 29835 14929 29838
rect 15700 29873 16110 30247
rect 19518 30317 19920 30320
rect 19518 30233 19523 30317
rect 19915 30233 19920 30317
rect 19518 30230 19920 30233
rect 19662 30056 19712 30059
rect 19662 30045 19665 30056
rect 16233 30042 19665 30045
rect 16233 29998 16236 30042
rect 16280 29998 19665 30042
rect 19709 29998 19712 30056
rect 16233 29995 19712 29998
rect 19726 29992 19776 29995
rect 19726 29981 19729 29992
rect 16233 29978 19729 29981
rect 16233 29934 16236 29978
rect 16280 29934 19729 29978
rect 19773 29934 19776 29992
rect 16233 29931 19776 29934
rect 15700 29847 15703 29873
rect 16107 29847 16110 29873
rect 5138 29818 5349 29821
rect 5138 29760 5141 29818
rect 5167 29760 5320 29818
rect 5346 29760 5349 29818
rect 5138 29757 5349 29760
rect 14611 29818 14822 29821
rect 14611 29760 14614 29818
rect 14640 29760 14793 29818
rect 14819 29760 14822 29818
rect 14611 29757 14822 29760
rect 4989 29587 5190 29590
rect 4989 29535 4992 29587
rect 5044 29535 5190 29587
rect 4989 29532 5190 29535
rect 14770 29587 14971 29590
rect 14770 29535 14916 29587
rect 14968 29535 14971 29587
rect 14770 29532 14971 29535
rect 40 29259 3060 29262
rect 40 29215 2863 29259
rect 3055 29215 3060 29259
rect 40 29212 3060 29215
rect 3677 29242 3727 29245
rect 3677 29198 3680 29242
rect 3724 29198 3727 29242
rect 3677 29195 3727 29198
rect 3677 29178 3727 29181
rect 3677 29134 3680 29178
rect 3724 29134 3727 29178
rect 3677 29131 3727 29134
rect 3850 29047 3853 29473
rect 4257 29047 4260 29473
rect 5031 29496 5242 29499
rect 5031 29438 5034 29496
rect 5060 29438 5213 29496
rect 5239 29438 5242 29496
rect 5031 29435 5242 29438
rect 14718 29496 14929 29499
rect 14718 29438 14721 29496
rect 14747 29438 14900 29496
rect 14926 29438 14929 29496
rect 14718 29435 14929 29438
rect 15700 29473 16110 29847
rect 16233 29642 16283 29645
rect 16233 29598 16236 29642
rect 16280 29598 16283 29642
rect 16233 29595 16283 29598
rect 16233 29578 16283 29581
rect 16233 29534 16236 29578
rect 16280 29534 16283 29578
rect 16233 29531 16283 29534
rect 4989 29187 5190 29190
rect 4989 29135 4992 29187
rect 5044 29135 5190 29187
rect 4989 29132 5190 29135
rect 14770 29187 14971 29190
rect 14770 29135 14916 29187
rect 14968 29135 14971 29187
rect 14770 29132 14971 29135
rect 3850 29042 4260 29047
rect 5031 29096 5242 29099
rect 5031 29038 5034 29096
rect 5060 29038 5213 29096
rect 5239 29038 5242 29096
rect 5031 29035 5242 29038
rect 14718 29096 14929 29099
rect 14718 29038 14721 29096
rect 14747 29038 14900 29096
rect 14926 29038 14929 29096
rect 15700 29047 15703 29473
rect 16107 29047 16110 29473
rect 40060 29262 40160 30712
rect 16233 29242 16283 29245
rect 16233 29198 16236 29242
rect 16280 29198 16283 29242
rect 39960 29212 40160 29262
rect 16233 29195 16283 29198
rect 16233 29178 16283 29181
rect 16233 29134 16236 29178
rect 16280 29134 16283 29178
rect 16233 29131 16283 29134
rect 15700 29042 16110 29047
rect 14718 29035 14929 29038
rect 40 29007 2730 29010
rect 40 28960 2683 29007
rect 2680 28949 2683 28960
rect 2727 28949 2730 29007
rect 17230 29007 19920 29010
rect 2680 28946 2730 28949
rect 5170 28998 5820 29000
rect 40 28917 2666 28920
rect 40 28870 2619 28917
rect 2616 28859 2619 28870
rect 2663 28859 2666 28917
rect 5170 28908 5175 28998
rect 5815 28908 5820 28998
rect 5170 28903 5820 28908
rect 14140 28998 14790 29003
rect 14140 28908 14145 28998
rect 14785 28908 14790 28998
rect 17230 28949 17233 29007
rect 17277 28960 19920 29007
rect 17277 28949 17280 28960
rect 17230 28946 17280 28949
rect 14140 28903 14790 28908
rect 17294 28917 19920 28920
rect 2616 28856 2666 28859
rect 17294 28859 17297 28917
rect 17341 28870 19920 28917
rect 17341 28859 17344 28870
rect 17294 28856 17344 28859
rect 40 28817 440 28820
rect 40 28733 43 28817
rect 435 28733 440 28817
rect 40 28730 440 28733
rect 19518 28817 19920 28820
rect 19518 28733 19523 28817
rect 19915 28733 19920 28817
rect 19518 28730 19920 28733
rect 40060 27762 40160 29212
rect 40 27759 3060 27762
rect 40 27715 2863 27759
rect 3055 27715 3060 27759
rect 40 27712 3060 27715
rect 39960 27712 40160 27762
rect 40 27507 2602 27510
rect 40 27460 2555 27507
rect 2552 27449 2555 27460
rect 2599 27449 2602 27507
rect 2552 27446 2602 27449
rect 17358 27507 19920 27510
rect 17358 27449 17361 27507
rect 17405 27460 19920 27507
rect 17405 27449 17408 27460
rect 17358 27446 17408 27449
rect 40 27417 2538 27420
rect 40 27370 2491 27417
rect 2488 27359 2491 27370
rect 2535 27359 2538 27417
rect 2488 27356 2538 27359
rect 17422 27417 19920 27420
rect 17422 27359 17425 27417
rect 17469 27370 19920 27417
rect 17469 27359 17472 27370
rect 17422 27356 17472 27359
rect 40 27317 440 27320
rect 40 27233 43 27317
rect 435 27233 440 27317
rect 40 27230 440 27233
rect 19518 27317 19920 27320
rect 19518 27233 19523 27317
rect 19915 27233 19920 27317
rect 19518 27230 19920 27233
rect 40060 26262 40160 27712
rect 40 26259 3060 26262
rect 40 26215 2863 26259
rect 3055 26215 3060 26259
rect 40 26212 3060 26215
rect 39960 26212 40160 26262
rect 40 26007 2474 26010
rect 40 25960 2427 26007
rect 2424 25949 2427 25960
rect 2471 25949 2474 26007
rect 2424 25946 2474 25949
rect 17486 26007 19920 26010
rect 17486 25949 17489 26007
rect 17533 25960 19920 26007
rect 17533 25949 17536 25960
rect 17486 25946 17536 25949
rect 40 25917 2410 25920
rect 40 25870 2363 25917
rect 2360 25859 2363 25870
rect 2407 25859 2410 25917
rect 2360 25856 2410 25859
rect 17550 25917 19920 25920
rect 17550 25859 17553 25917
rect 17597 25870 19920 25917
rect 17597 25859 17600 25870
rect 17550 25856 17600 25859
rect 40 25817 440 25820
rect 40 25733 43 25817
rect 435 25733 440 25817
rect 40 25730 440 25733
rect 19518 25817 19920 25820
rect 19518 25733 19523 25817
rect 19915 25733 19920 25817
rect 19518 25730 19920 25733
rect 40060 24762 40160 26212
rect 40 24759 3060 24762
rect 40 24715 2863 24759
rect 3055 24715 3060 24759
rect 40 24712 3060 24715
rect 39960 24712 40160 24762
rect 40 24507 2346 24510
rect 40 24460 2299 24507
rect 2296 24449 2299 24460
rect 2343 24449 2346 24507
rect 2296 24446 2346 24449
rect 17614 24507 19920 24510
rect 17614 24449 17617 24507
rect 17661 24460 19920 24507
rect 17661 24449 17664 24460
rect 17614 24446 17664 24449
rect 40 24417 2282 24420
rect 40 24370 2235 24417
rect 2232 24359 2235 24370
rect 2279 24359 2282 24417
rect 2232 24356 2282 24359
rect 17678 24417 19920 24420
rect 17678 24359 17681 24417
rect 17725 24370 19920 24417
rect 17725 24359 17728 24370
rect 17678 24356 17728 24359
rect 40 24317 440 24320
rect 40 24233 43 24317
rect 435 24233 440 24317
rect 40 24230 440 24233
rect 19518 24317 19920 24320
rect 19518 24233 19523 24317
rect 19915 24233 19920 24317
rect 19518 24230 19920 24233
rect 40060 23262 40160 24712
rect 40 23259 3060 23262
rect 40 23215 2863 23259
rect 3055 23215 3060 23259
rect 40 23212 3060 23215
rect 39960 23212 40160 23262
rect 40 23007 2218 23010
rect 40 22960 2171 23007
rect 2168 22949 2171 22960
rect 2215 22949 2218 23007
rect 2168 22946 2218 22949
rect 17742 23007 19920 23010
rect 17742 22949 17745 23007
rect 17789 22960 19920 23007
rect 17789 22949 17792 22960
rect 17742 22946 17792 22949
rect 40 22917 2154 22920
rect 40 22870 2107 22917
rect 2104 22859 2107 22870
rect 2151 22859 2154 22917
rect 2104 22856 2154 22859
rect 17806 22917 19920 22920
rect 17806 22859 17809 22917
rect 17853 22870 19920 22917
rect 17853 22859 17856 22870
rect 17806 22856 17856 22859
rect 40 22817 440 22820
rect 40 22733 43 22817
rect 435 22733 440 22817
rect 40 22730 440 22733
rect 19518 22817 19920 22820
rect 19518 22733 19523 22817
rect 19915 22733 19920 22817
rect 19518 22730 19920 22733
rect 40060 21762 40160 23212
rect 40 21759 3060 21762
rect 40 21715 2863 21759
rect 3055 21715 3060 21759
rect 40 21712 3060 21715
rect 39960 21712 40160 21762
rect 40 21507 2090 21510
rect 40 21460 2043 21507
rect 2040 21449 2043 21460
rect 2087 21449 2090 21507
rect 2040 21446 2090 21449
rect 17870 21507 19920 21510
rect 17870 21449 17873 21507
rect 17917 21460 19920 21507
rect 17917 21449 17920 21460
rect 17870 21446 17920 21449
rect 40 21417 2026 21420
rect 40 21370 1979 21417
rect 1976 21359 1979 21370
rect 2023 21359 2026 21417
rect 1976 21356 2026 21359
rect 17934 21417 19920 21420
rect 17934 21359 17937 21417
rect 17981 21370 19920 21417
rect 17981 21359 17984 21370
rect 17934 21356 17984 21359
rect 40 21317 440 21320
rect 40 21233 43 21317
rect 435 21233 440 21317
rect 19518 21317 19920 21320
rect 40 21230 440 21233
rect 5170 21295 5820 21300
rect 5170 21105 5175 21295
rect 5815 21105 5820 21295
rect 5170 21100 5820 21105
rect 14140 21295 14790 21300
rect 14140 21105 14145 21295
rect 14785 21105 14790 21295
rect 19518 21233 19523 21317
rect 19915 21233 19920 21317
rect 19518 21230 19920 21233
rect 14140 21100 14790 21105
rect 40060 20262 40160 21712
rect 40 20259 3060 20262
rect 40 20215 2863 20259
rect 3055 20215 3060 20259
rect 40 20212 3060 20215
rect 39960 20212 40160 20262
rect 40 20007 1962 20010
rect 40 19960 1915 20007
rect 1912 19949 1915 19960
rect 1959 19949 1962 20007
rect 1912 19946 1962 19949
rect 17998 20007 19920 20010
rect 17998 19949 18001 20007
rect 18045 19960 19920 20007
rect 18045 19949 18048 19960
rect 17998 19946 18048 19949
rect 40 19917 1898 19920
rect 40 19870 1851 19917
rect 1848 19859 1851 19870
rect 1895 19859 1898 19917
rect 18062 19917 19920 19920
rect 1848 19856 1898 19859
rect 40 19817 440 19820
rect 40 19780 43 19817
rect 38 19563 43 19780
rect 435 19780 440 19817
rect 3857 19780 3884 19900
rect 15957 19780 15984 19900
rect 18062 19859 18065 19917
rect 18109 19870 19920 19917
rect 18109 19859 18112 19870
rect 18062 19856 18112 19859
rect 19518 19817 19920 19820
rect 19518 19780 19523 19817
rect 435 19563 19523 19780
rect 19915 19563 19920 19817
rect 38 19560 19920 19563
rect 38 19558 440 19560
rect 10430 19277 10650 19560
rect 10965 19460 11095 19465
rect 10965 19340 10970 19460
rect 11090 19340 11095 19460
rect 10965 19335 11095 19340
rect 10430 19066 10593 19277
rect 10646 19066 10650 19277
rect 10430 19060 10650 19066
rect 10999 19270 11040 19335
rect 10999 19060 11002 19270
rect 11037 19060 11040 19270
rect 10999 19057 11040 19060
rect 11114 19273 11174 19276
rect 11114 19063 11117 19273
rect 11171 19063 11174 19273
rect 40 18759 3060 18762
rect 40 18715 2863 18759
rect 3055 18715 3060 18759
rect 40 18712 3060 18715
rect 40 18507 1834 18510
rect 40 18460 1787 18507
rect 1784 18449 1787 18460
rect 1831 18449 1834 18507
rect 1784 18446 1834 18449
rect 40 18417 1770 18420
rect 40 18370 1723 18417
rect 1720 18359 1723 18370
rect 1767 18359 1770 18417
rect 11114 18375 11174 19063
rect 40060 18762 40160 20212
rect 39960 18712 40160 18762
rect 18126 18507 19920 18510
rect 18126 18449 18129 18507
rect 18173 18460 19920 18507
rect 18173 18449 18176 18460
rect 18126 18446 18176 18449
rect 18190 18417 19920 18420
rect 1720 18356 1770 18359
rect 11065 18370 11195 18375
rect 40 18317 440 18320
rect 40 18233 43 18317
rect 435 18233 440 18317
rect 11065 18250 11070 18370
rect 11190 18250 11195 18370
rect 18190 18359 18193 18417
rect 18237 18370 19920 18417
rect 18237 18359 18240 18370
rect 18190 18356 18240 18359
rect 11065 18245 11195 18250
rect 19518 18317 19920 18320
rect 40 18230 440 18233
rect 19518 18233 19523 18317
rect 19915 18233 19920 18317
rect 19518 18230 19920 18233
rect 40060 17262 40160 18712
rect 40 17259 3060 17262
rect 40 17215 2863 17259
rect 3055 17215 3060 17259
rect 40 17212 3060 17215
rect 39960 17212 40160 17262
rect 40 17007 1706 17010
rect 40 16960 1659 17007
rect 1656 16949 1659 16960
rect 1703 16949 1706 17007
rect 1656 16946 1706 16949
rect 18254 17007 19920 17010
rect 18254 16949 18257 17007
rect 18301 16960 19920 17007
rect 18301 16949 18304 16960
rect 18254 16946 18304 16949
rect 40 16917 1642 16920
rect 40 16870 1595 16917
rect 1592 16859 1595 16870
rect 1639 16859 1642 16917
rect 1592 16856 1642 16859
rect 18318 16917 19920 16920
rect 18318 16859 18321 16917
rect 18365 16870 19920 16917
rect 18365 16859 18368 16870
rect 18318 16856 18368 16859
rect 40 16817 440 16820
rect 40 16733 43 16817
rect 435 16733 440 16817
rect 40 16730 440 16733
rect 19518 16817 19920 16820
rect 19518 16733 19523 16817
rect 19915 16733 19920 16817
rect 19518 16730 19920 16733
rect 40060 15762 40160 17212
rect 40 15759 3060 15762
rect 40 15715 2863 15759
rect 3055 15715 3060 15759
rect 40 15712 3060 15715
rect 39960 15712 40160 15762
rect 40 15507 1578 15510
rect 40 15460 1531 15507
rect 1528 15449 1531 15460
rect 1575 15449 1578 15507
rect 1528 15446 1578 15449
rect 18382 15507 19920 15510
rect 18382 15449 18385 15507
rect 18429 15460 19920 15507
rect 18429 15449 18432 15460
rect 18382 15446 18432 15449
rect 40 15417 1514 15420
rect 40 15370 1467 15417
rect 1464 15359 1467 15370
rect 1511 15359 1514 15417
rect 1464 15356 1514 15359
rect 18446 15417 19920 15420
rect 18446 15359 18449 15417
rect 18493 15370 19920 15417
rect 18493 15359 18496 15370
rect 18446 15356 18496 15359
rect 40 15317 440 15320
rect 40 15233 43 15317
rect 435 15233 440 15317
rect 40 15230 440 15233
rect 19518 15317 19920 15320
rect 19518 15233 19523 15317
rect 19915 15233 19920 15317
rect 19518 15230 19920 15233
rect 40060 14262 40160 15712
rect 40 14259 3060 14262
rect 40 14215 2863 14259
rect 3055 14215 3060 14259
rect 40 14212 3060 14215
rect 39960 14212 40160 14262
rect 40 14007 1450 14010
rect 40 13960 1403 14007
rect 1400 13949 1403 13960
rect 1447 13949 1450 14007
rect 1400 13946 1450 13949
rect 18510 14007 19920 14010
rect 18510 13949 18513 14007
rect 18557 13960 19920 14007
rect 18557 13949 18560 13960
rect 18510 13946 18560 13949
rect 40 13917 1386 13920
rect 40 13870 1339 13917
rect 1336 13859 1339 13870
rect 1383 13859 1386 13917
rect 1336 13856 1386 13859
rect 18574 13917 19920 13920
rect 18574 13859 18577 13917
rect 18621 13870 19920 13917
rect 18621 13859 18624 13870
rect 18574 13856 18624 13859
rect 40 13817 440 13820
rect 40 13733 43 13817
rect 435 13733 440 13817
rect 40 13730 440 13733
rect 19518 13817 19920 13820
rect 19518 13733 19523 13817
rect 19915 13733 19920 13817
rect 19518 13730 19920 13733
rect 40060 12762 40160 14212
rect 40 12759 3060 12762
rect 40 12715 2863 12759
rect 3055 12715 3060 12759
rect 40 12712 3060 12715
rect 39960 12712 40160 12762
rect 40 12507 1322 12510
rect 40 12460 1275 12507
rect 1272 12449 1275 12460
rect 1319 12449 1322 12507
rect 1272 12446 1322 12449
rect 18638 12507 19920 12510
rect 18638 12449 18641 12507
rect 18685 12460 19920 12507
rect 18685 12449 18688 12460
rect 18638 12446 18688 12449
rect 40 12417 1258 12420
rect 40 12370 1211 12417
rect 1208 12359 1211 12370
rect 1255 12359 1258 12417
rect 1208 12356 1258 12359
rect 18702 12417 19920 12420
rect 18702 12359 18705 12417
rect 18749 12370 19920 12417
rect 18749 12359 18752 12370
rect 18702 12356 18752 12359
rect 40 12317 440 12320
rect 40 12233 43 12317
rect 435 12233 440 12317
rect 40 12230 440 12233
rect 19518 12317 19920 12320
rect 19518 12233 19523 12317
rect 19915 12233 19920 12317
rect 19518 12230 19920 12233
rect 40060 11262 40160 12712
rect 40 11259 3060 11262
rect 40 11215 2863 11259
rect 3055 11215 3060 11259
rect 40 11212 3060 11215
rect 39960 11212 40160 11262
rect 40 11007 1194 11010
rect 40 10960 1147 11007
rect 1144 10949 1147 10960
rect 1191 10949 1194 11007
rect 1144 10946 1194 10949
rect 18766 11007 19920 11010
rect 18766 10949 18769 11007
rect 18813 10960 19920 11007
rect 18813 10949 18816 10960
rect 18766 10946 18816 10949
rect 40 10917 1130 10920
rect 40 10870 1083 10917
rect 1080 10859 1083 10870
rect 1127 10859 1130 10917
rect 1080 10856 1130 10859
rect 18830 10917 19920 10920
rect 18830 10859 18833 10917
rect 18877 10870 19920 10917
rect 18877 10859 18880 10870
rect 18830 10856 18880 10859
rect 40 10817 440 10820
rect 40 10733 43 10817
rect 435 10733 440 10817
rect 40 10730 440 10733
rect 19518 10817 19920 10820
rect 19518 10733 19523 10817
rect 19915 10733 19920 10817
rect 19518 10730 19920 10733
rect 40060 9762 40160 11212
rect 40 9759 3060 9762
rect 40 9715 2863 9759
rect 3055 9715 3060 9759
rect 40 9712 3060 9715
rect 39960 9712 40160 9762
rect 40 9507 1066 9510
rect 40 9460 1019 9507
rect 1016 9449 1019 9460
rect 1063 9449 1066 9507
rect 1016 9446 1066 9449
rect 18894 9507 19920 9510
rect 18894 9449 18897 9507
rect 18941 9460 19920 9507
rect 18941 9449 18944 9460
rect 18894 9446 18944 9449
rect 40 9417 1002 9420
rect 40 9370 955 9417
rect 952 9359 955 9370
rect 999 9359 1002 9417
rect 952 9356 1002 9359
rect 18958 9417 19920 9420
rect 18958 9359 18961 9417
rect 19005 9370 19920 9417
rect 19005 9359 19008 9370
rect 18958 9356 19008 9359
rect 40 9317 440 9320
rect 40 9233 43 9317
rect 435 9233 440 9317
rect 40 9230 440 9233
rect 19518 9317 19920 9320
rect 19518 9233 19523 9317
rect 19915 9233 19920 9317
rect 19518 9230 19920 9233
rect 40060 8262 40160 9712
rect 40 8259 3060 8262
rect 40 8215 2863 8259
rect 3055 8215 3060 8259
rect 40 8212 3060 8215
rect 39960 8212 40160 8262
rect 40 8007 938 8010
rect 40 7960 891 8007
rect 888 7949 891 7960
rect 935 7949 938 8007
rect 888 7946 938 7949
rect 19022 8007 19920 8010
rect 19022 7949 19025 8007
rect 19069 7960 19920 8007
rect 19069 7949 19072 7960
rect 19022 7946 19072 7949
rect 40 7917 874 7920
rect 40 7870 827 7917
rect 824 7859 827 7870
rect 871 7859 874 7917
rect 824 7856 874 7859
rect 19086 7917 19920 7920
rect 19086 7859 19089 7917
rect 19133 7870 19920 7917
rect 19133 7859 19136 7870
rect 19086 7856 19136 7859
rect 40 7817 440 7820
rect 40 7733 43 7817
rect 435 7733 440 7817
rect 40 7730 440 7733
rect 19518 7817 19920 7820
rect 19518 7733 19523 7817
rect 19915 7733 19920 7817
rect 19518 7730 19920 7733
rect 40060 6762 40160 8212
rect 40 6759 3060 6762
rect 40 6715 2863 6759
rect 3055 6715 3060 6759
rect 40 6712 3060 6715
rect 39960 6712 40160 6762
rect 40 6507 810 6510
rect 40 6460 763 6507
rect 760 6449 763 6460
rect 807 6449 810 6507
rect 760 6446 810 6449
rect 19150 6507 19920 6510
rect 19150 6449 19153 6507
rect 19197 6460 19920 6507
rect 19197 6449 19200 6460
rect 19150 6446 19200 6449
rect 40 6417 746 6420
rect 40 6370 699 6417
rect 696 6359 699 6370
rect 743 6359 746 6417
rect 696 6356 746 6359
rect 19214 6417 19920 6420
rect 19214 6359 19217 6417
rect 19261 6370 19920 6417
rect 19261 6359 19264 6370
rect 19214 6356 19264 6359
rect 40 6317 440 6320
rect 40 6233 43 6317
rect 435 6233 440 6317
rect 40 6230 440 6233
rect 19518 6317 19920 6320
rect 19518 6233 19523 6317
rect 19915 6233 19920 6317
rect 19518 6230 19920 6233
rect 8774 6201 12968 6204
rect 8774 6199 12871 6201
rect 8774 6109 8779 6199
rect 8969 6109 12871 6199
rect 8774 6107 12871 6109
rect 12965 6107 12968 6201
rect 8774 6104 12968 6107
rect 9042 6033 13106 6036
rect 9042 6031 13009 6033
rect 9042 5941 9047 6031
rect 9237 5941 13009 6031
rect 9042 5939 13009 5941
rect 13103 5939 13106 6033
rect 9042 5936 13106 5939
rect 9310 5865 13244 5868
rect 9310 5863 13147 5865
rect 9310 5773 9315 5863
rect 9505 5773 13147 5863
rect 9310 5771 13147 5773
rect 13241 5771 13244 5865
rect 9310 5768 13244 5771
rect 9578 5697 13382 5700
rect 9578 5695 13285 5697
rect 9578 5605 9583 5695
rect 9773 5605 13285 5695
rect 9578 5603 13285 5605
rect 13379 5603 13382 5697
rect 9578 5600 13382 5603
rect 12868 5577 12968 5580
rect 12868 5483 12871 5577
rect 12965 5483 12968 5577
rect 12868 5480 12968 5483
rect 13006 5577 13106 5580
rect 13006 5483 13009 5577
rect 13103 5483 13106 5577
rect 13006 5480 13106 5483
rect 13144 5577 13244 5580
rect 13144 5483 13147 5577
rect 13241 5483 13244 5577
rect 13144 5480 13244 5483
rect 40060 5262 40160 6712
rect 40 5259 3060 5262
rect 40 5215 2863 5259
rect 3055 5215 3060 5259
rect 40 5212 3060 5215
rect 39960 5212 40160 5262
rect 40 5007 682 5010
rect 40 4960 635 5007
rect 632 4949 635 4960
rect 679 4949 682 5007
rect 632 4946 682 4949
rect 19278 5007 19920 5010
rect 19278 4949 19281 5007
rect 19325 4960 19920 5007
rect 19325 4949 19328 4960
rect 19278 4946 19328 4949
rect 40 4917 618 4920
rect 40 4870 571 4917
rect 568 4859 571 4870
rect 615 4859 618 4917
rect 568 4856 618 4859
rect 19342 4917 19920 4920
rect 19342 4859 19345 4917
rect 19389 4870 19920 4917
rect 19389 4859 19392 4870
rect 19342 4856 19392 4859
rect 40 4817 440 4820
rect 40 4733 43 4817
rect 435 4733 440 4817
rect 40 4730 440 4733
rect 19518 4817 19920 4820
rect 19518 4733 19523 4817
rect 19915 4733 19920 4817
rect 19518 4730 19920 4733
rect 40060 3762 40160 5212
rect 40 3759 3060 3762
rect 40 3715 2863 3759
rect 3055 3715 3060 3759
rect 40 3712 3060 3715
rect 39960 3712 40160 3762
rect 40 3507 554 3510
rect 40 3460 507 3507
rect 504 3449 507 3460
rect 551 3449 554 3507
rect 504 3446 554 3449
rect 19406 3507 19920 3510
rect 19406 3449 19409 3507
rect 19453 3460 19920 3507
rect 19453 3449 19456 3460
rect 19406 3446 19456 3449
rect 40 3417 490 3420
rect 40 3370 443 3417
rect 440 3359 443 3370
rect 487 3359 490 3417
rect 440 3356 490 3359
rect 19470 3417 19920 3420
rect 19470 3359 19473 3417
rect 19517 3370 19920 3417
rect 19517 3359 19520 3370
rect 19470 3356 19520 3359
rect 40 3317 440 3320
rect 40 3233 43 3317
rect 435 3233 440 3317
rect 40 3230 440 3233
rect 19518 3317 19920 3320
rect 19518 3233 19523 3317
rect 19915 3233 19920 3317
rect 19518 3230 19920 3233
rect 12700 2625 15100 2630
rect 40 2259 3060 2262
rect 40 2215 2863 2259
rect 3055 2215 3060 2259
rect 40 2212 3060 2215
rect 6811 2156 6869 2159
rect 6811 2130 6814 2156
rect 6866 2130 6869 2156
rect 6083 2049 6141 2052
rect 6083 2023 6086 2049
rect 6138 2023 6141 2049
rect 40 2007 426 2010
rect 40 1960 379 2007
rect 376 1949 379 1960
rect 423 1949 426 2007
rect 376 1946 426 1949
rect 40 1917 362 1920
rect 40 1870 315 1917
rect 312 1859 315 1870
rect 359 1859 362 1917
rect 312 1856 362 1859
rect 6083 1870 6141 2023
rect 6483 2049 6541 2052
rect 6483 2023 6486 2049
rect 6538 2023 6541 2049
rect 6083 1844 6086 1870
rect 6138 1844 6141 1870
rect 6083 1841 6141 1844
rect 6180 1854 6238 2000
rect 40 1817 440 1820
rect 40 1733 43 1817
rect 435 1733 440 1817
rect 6180 1802 6183 1854
rect 6235 1802 6238 1854
rect 6483 1870 6541 2023
rect 6483 1844 6486 1870
rect 6538 1844 6541 1870
rect 6483 1841 6541 1844
rect 6580 1854 6638 2000
rect 6811 1977 6869 2130
rect 7611 2156 7669 2159
rect 7611 2130 7614 2156
rect 7666 2130 7669 2156
rect 6811 1951 6814 1977
rect 6866 1951 6869 1977
rect 6811 1948 6869 1951
rect 6883 2049 6941 2052
rect 6883 2023 6886 2049
rect 6938 2023 6941 2049
rect 6180 1799 6238 1802
rect 6580 1802 6583 1854
rect 6635 1802 6638 1854
rect 6883 1870 6941 2023
rect 7283 2049 7341 2052
rect 7283 2023 7286 2049
rect 7338 2023 7341 2049
rect 6883 1844 6886 1870
rect 6938 1844 6941 1870
rect 6883 1841 6941 1844
rect 6980 1854 7038 2000
rect 6580 1799 6638 1802
rect 6980 1802 6983 1854
rect 7035 1802 7038 1854
rect 7283 1870 7341 2023
rect 7283 1844 7286 1870
rect 7338 1844 7341 1870
rect 7283 1841 7341 1844
rect 7380 1854 7438 2000
rect 7611 1977 7669 2130
rect 8411 2156 8469 2159
rect 8411 2130 8414 2156
rect 8466 2130 8469 2156
rect 7611 1951 7614 1977
rect 7666 1951 7669 1977
rect 7611 1948 7669 1951
rect 7683 2049 7741 2052
rect 7683 2023 7686 2049
rect 7738 2023 7741 2049
rect 6980 1799 7038 1802
rect 7380 1802 7383 1854
rect 7435 1802 7438 1854
rect 7683 1870 7741 2023
rect 8083 2049 8141 2052
rect 8083 2023 8086 2049
rect 8138 2023 8141 2049
rect 7683 1844 7686 1870
rect 7738 1844 7741 1870
rect 7683 1841 7741 1844
rect 7780 1854 7838 2000
rect 7380 1799 7438 1802
rect 7780 1802 7783 1854
rect 7835 1802 7838 1854
rect 8083 1870 8141 2023
rect 8083 1844 8086 1870
rect 8138 1844 8141 1870
rect 8083 1841 8141 1844
rect 8180 1854 8238 2000
rect 8411 1977 8469 2130
rect 9211 2156 9269 2159
rect 9211 2130 9214 2156
rect 9266 2130 9269 2156
rect 8411 1951 8414 1977
rect 8466 1951 8469 1977
rect 8411 1948 8469 1951
rect 8483 2049 8541 2052
rect 8483 2023 8486 2049
rect 8538 2023 8541 2049
rect 7780 1799 7838 1802
rect 8180 1802 8183 1854
rect 8235 1802 8238 1854
rect 8483 1870 8541 2023
rect 8883 2049 8941 2052
rect 8883 2023 8886 2049
rect 8938 2023 8941 2049
rect 8483 1844 8486 1870
rect 8538 1844 8541 1870
rect 8483 1841 8541 1844
rect 8580 1854 8638 2000
rect 8180 1799 8238 1802
rect 8580 1802 8583 1854
rect 8635 1802 8638 1854
rect 8883 1870 8941 2023
rect 8883 1844 8886 1870
rect 8938 1844 8941 1870
rect 8883 1841 8941 1844
rect 8980 1854 9038 2000
rect 9211 1977 9269 2130
rect 10011 2156 10069 2159
rect 10011 2130 10014 2156
rect 10066 2130 10069 2156
rect 9211 1951 9214 1977
rect 9266 1951 9269 1977
rect 9211 1948 9269 1951
rect 9283 2049 9341 2052
rect 9283 2023 9286 2049
rect 9338 2023 9341 2049
rect 8580 1799 8638 1802
rect 8980 1802 8983 1854
rect 9035 1802 9038 1854
rect 9283 1870 9341 2023
rect 9683 2049 9741 2052
rect 9683 2023 9686 2049
rect 9738 2023 9741 2049
rect 9283 1844 9286 1870
rect 9338 1844 9341 1870
rect 9283 1841 9341 1844
rect 9380 1854 9438 2000
rect 8980 1799 9038 1802
rect 9380 1802 9383 1854
rect 9435 1802 9438 1854
rect 9683 1870 9741 2023
rect 9683 1844 9686 1870
rect 9738 1844 9741 1870
rect 9683 1841 9741 1844
rect 9780 1854 9838 2000
rect 10011 1977 10069 2130
rect 10811 2156 10869 2159
rect 10811 2130 10814 2156
rect 10866 2130 10869 2156
rect 10011 1951 10014 1977
rect 10066 1951 10069 1977
rect 10011 1948 10069 1951
rect 10083 2049 10141 2052
rect 10083 2023 10086 2049
rect 10138 2023 10141 2049
rect 9380 1799 9438 1802
rect 9780 1802 9783 1854
rect 9835 1802 9838 1854
rect 10083 1870 10141 2023
rect 10483 2049 10541 2052
rect 10483 2023 10486 2049
rect 10538 2023 10541 2049
rect 10083 1844 10086 1870
rect 10138 1844 10141 1870
rect 10083 1841 10141 1844
rect 10180 1854 10238 2000
rect 9780 1799 9838 1802
rect 10180 1802 10183 1854
rect 10235 1802 10238 1854
rect 10483 1870 10541 2023
rect 10483 1844 10486 1870
rect 10538 1844 10541 1870
rect 10483 1841 10541 1844
rect 10580 1854 10638 2000
rect 10811 1977 10869 2130
rect 11611 2156 11669 2159
rect 11611 2130 11614 2156
rect 11666 2130 11669 2156
rect 12700 2135 14903 2625
rect 15097 2135 15100 2625
rect 40060 2262 40160 3712
rect 39960 2212 40160 2262
rect 12700 2130 15100 2135
rect 10811 1951 10814 1977
rect 10866 1951 10869 1977
rect 10811 1948 10869 1951
rect 10883 2049 10941 2052
rect 10883 2023 10886 2049
rect 10938 2023 10941 2049
rect 10180 1799 10238 1802
rect 10580 1802 10583 1854
rect 10635 1802 10638 1854
rect 10883 1870 10941 2023
rect 11283 2049 11341 2052
rect 11283 2023 11286 2049
rect 11338 2023 11341 2049
rect 10883 1844 10886 1870
rect 10938 1844 10941 1870
rect 10883 1841 10941 1844
rect 10980 1854 11038 2000
rect 10580 1799 10638 1802
rect 10980 1802 10983 1854
rect 11035 1802 11038 1854
rect 11283 1870 11341 2023
rect 11283 1844 11286 1870
rect 11338 1844 11341 1870
rect 11283 1841 11341 1844
rect 11380 1854 11438 2000
rect 11611 1977 11669 2130
rect 12430 2080 12530 2130
rect 12430 2075 14340 2080
rect 11611 1951 11614 1977
rect 11666 1951 11669 1977
rect 11611 1948 11669 1951
rect 11683 2049 11741 2052
rect 11683 2023 11686 2049
rect 11738 2023 11741 2049
rect 10980 1799 11038 1802
rect 11380 1802 11383 1854
rect 11435 1802 11438 1854
rect 11683 1870 11741 2023
rect 12083 2049 12141 2052
rect 12083 2023 12086 2049
rect 12138 2023 12141 2049
rect 11683 1844 11686 1870
rect 11738 1844 11741 1870
rect 11683 1841 11741 1844
rect 11780 1854 11838 2000
rect 11380 1799 11438 1802
rect 11780 1802 11783 1854
rect 11835 1802 11838 1854
rect 12083 1870 12141 2023
rect 12083 1844 12086 1870
rect 12138 1844 12141 1870
rect 12083 1841 12141 1844
rect 12180 1854 12238 2000
rect 11780 1799 11838 1802
rect 12180 1802 12183 1854
rect 12235 1802 12238 1854
rect 12180 1799 12238 1802
rect 12430 1977 14143 2075
rect 12430 1903 12443 1977
rect 12517 1903 14143 1977
rect 40 1730 440 1733
rect 12430 1585 14143 1903
rect 14337 1585 14340 2075
rect 19534 2007 19920 2010
rect 19534 1949 19537 2007
rect 19581 1960 19920 2007
rect 19581 1949 19584 1960
rect 19534 1946 19584 1949
rect 19598 1917 19920 1920
rect 19598 1859 19601 1917
rect 19645 1870 19920 1917
rect 19645 1859 19648 1870
rect 19598 1856 19648 1859
rect 19518 1817 19920 1820
rect 19518 1733 19523 1817
rect 19915 1733 19920 1817
rect 19518 1730 19920 1733
rect 12430 1580 14340 1585
rect 6080 987 16330 990
rect 40 759 3060 762
rect 40 715 2863 759
rect 3055 715 3060 759
rect 40 712 3060 715
rect 6080 593 6090 987
rect 6116 593 6490 987
rect 6516 593 6890 987
rect 6916 593 7290 987
rect 7316 593 7690 987
rect 7716 593 8090 987
rect 8116 593 8490 987
rect 8516 593 8890 987
rect 8916 593 9290 987
rect 9316 593 9690 987
rect 9716 593 10090 987
rect 10116 593 10490 987
rect 10516 593 10890 987
rect 10916 593 11290 987
rect 11316 593 11690 987
rect 11716 593 12090 987
rect 12116 985 16330 987
rect 12116 595 15675 985
rect 16325 595 16330 985
rect 40060 849 40160 2212
rect 40060 832 40242 849
rect 40060 762 40100 832
rect 39960 712 40100 762
rect 40220 712 40242 832
rect 40093 705 40242 712
rect 12116 593 16330 595
rect 6080 590 16330 593
rect 40 507 298 510
rect 40 460 251 507
rect 248 449 251 460
rect 295 449 298 507
rect 248 446 298 449
rect 19662 507 19920 510
rect 19662 449 19665 507
rect 19709 460 19920 507
rect 19709 449 19712 460
rect 19662 446 19712 449
rect 40 417 234 420
rect 40 370 187 417
rect 184 359 187 370
rect 231 359 234 417
rect 184 356 234 359
rect 19726 417 19920 420
rect 19726 359 19729 417
rect 19773 370 19920 417
rect 19773 359 19776 370
rect 19726 356 19776 359
rect 40 317 440 320
rect 40 233 43 317
rect 435 280 440 317
rect 19518 317 19920 320
rect 435 277 1139 280
rect 435 233 1092 277
rect 1136 233 1139 277
rect 40 230 1139 233
rect 19518 233 19523 317
rect 19915 233 19920 317
rect 19518 230 19920 233
rect 7281 166 7479 169
rect 7281 140 7284 166
rect 7310 140 7450 166
rect 7476 140 7479 166
rect 7281 137 7479 140
rect 7027 120 7425 123
rect 7027 94 7030 120
rect 7056 94 7396 120
rect 7422 94 7425 120
rect 7027 91 7425 94
rect 6281 74 7879 77
rect 6281 48 6284 74
rect 6310 48 7850 74
rect 7876 48 7879 74
rect 6281 45 7879 48
rect 6027 28 7825 31
rect 6027 2 6030 28
rect 6056 2 7796 28
rect 7822 2 7825 28
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -220 -5 -140 0
rect 6027 -1 7825 2
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect 20100 -5 20180 0
rect 1281 -18 8279 -15
rect 1281 -44 1284 -18
rect 1310 -44 8250 -18
rect 8276 -44 8279 -18
rect 1281 -47 8279 -44
rect -220 -80 -140 -75
rect 1027 -64 8225 -61
rect 1027 -90 1030 -64
rect 1056 -90 8196 -64
rect 8222 -90 8225 -64
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
rect 1027 -93 8225 -90
rect -14 -110 19973 -107
rect -14 -136 -11 -110
rect 15 -136 12250 -110
rect 12276 -136 19944 -110
rect 19970 -136 19973 -110
rect -14 -139 19973 -136
rect -268 -156 20227 -153
rect -268 -182 -265 -156
rect -239 -182 12196 -156
rect 12222 -182 20198 -156
rect 20224 -182 20227 -156
rect -268 -185 20227 -182
rect -2016 -202 21975 -199
rect -2016 -228 -2011 -202
rect -1985 -228 11850 -202
rect 11876 -228 21944 -202
rect 21970 -228 21975 -202
rect -2016 -231 21975 -228
rect -2270 -248 22229 -245
rect -2270 -274 -2265 -248
rect -2239 -274 11796 -248
rect 11822 -274 22198 -248
rect 22224 -274 22229 -248
rect -2270 -277 22229 -274
rect -4016 -294 23975 -291
rect -4016 -320 -4011 -294
rect -3985 -320 11450 -294
rect 11476 -320 23944 -294
rect 23970 -320 23975 -294
rect -4016 -323 23975 -320
rect -4270 -340 24229 -337
rect -4270 -366 -4265 -340
rect -4239 -366 11396 -340
rect 11422 -366 24198 -340
rect 24224 -366 24229 -340
rect -4270 -369 24229 -366
rect -6016 -386 25975 -383
rect -6016 -412 -6011 -386
rect -5985 -412 11050 -386
rect 11076 -412 25944 -386
rect 25970 -412 25975 -386
rect -6016 -415 25975 -412
rect -6270 -432 26229 -429
rect -6270 -458 -6265 -432
rect -6239 -458 10996 -432
rect 11022 -458 26198 -432
rect 26224 -458 26229 -432
rect -6270 -461 26229 -458
rect -8016 -478 27975 -475
rect -8016 -504 -8011 -478
rect -7985 -504 10650 -478
rect 10676 -504 27944 -478
rect 27970 -504 27975 -478
rect -8016 -507 27975 -504
rect -8270 -524 28229 -521
rect -8270 -550 -8265 -524
rect -8239 -550 10596 -524
rect 10622 -550 28198 -524
rect 28224 -550 28229 -524
rect -8270 -553 28229 -550
rect -10016 -570 29975 -567
rect -10016 -596 -10011 -570
rect -9985 -596 10250 -570
rect 10276 -596 29944 -570
rect 29970 -596 29975 -570
rect -10016 -599 29975 -596
rect -10270 -616 30229 -613
rect -10270 -642 -10265 -616
rect -10239 -642 10196 -616
rect 10222 -642 30198 -616
rect 30224 -642 30229 -616
rect -10270 -645 30229 -642
rect -12016 -662 31975 -659
rect -12016 -688 -12011 -662
rect -11985 -688 9850 -662
rect 9876 -688 31944 -662
rect 31970 -688 31975 -662
rect -12016 -691 31975 -688
rect -12270 -708 32229 -705
rect -12270 -734 -12265 -708
rect -12239 -734 9796 -708
rect 9822 -734 32198 -708
rect 32224 -734 32229 -708
rect -12270 -737 32229 -734
rect -14016 -754 33975 -751
rect -14016 -780 -14011 -754
rect -13985 -780 9450 -754
rect 9476 -780 33944 -754
rect 33970 -780 33975 -754
rect -14016 -783 33975 -780
rect -14270 -800 34229 -797
rect -14270 -826 -14265 -800
rect -14239 -826 9396 -800
rect 9422 -826 34198 -800
rect 34224 -826 34229 -800
rect -14270 -829 34229 -826
rect -16014 -846 35973 -843
rect -16014 -872 -16011 -846
rect -15985 -872 9050 -846
rect 9076 -872 35944 -846
rect 35970 -872 35973 -846
rect -16014 -875 35973 -872
rect -16268 -892 36227 -889
rect -16268 -918 -16265 -892
rect -16239 -918 8996 -892
rect 9022 -918 36198 -892
rect 36224 -918 36227 -892
rect -16268 -921 36227 -918
rect -18014 -938 37973 -935
rect -18014 -964 -18011 -938
rect -17985 -964 8650 -938
rect 8676 -964 37944 -938
rect 37970 -964 37973 -938
rect -18014 -967 37973 -964
rect -18268 -984 38229 -981
rect -18268 -1010 -18265 -984
rect -18239 -1010 8596 -984
rect 8622 -1010 38198 -984
rect 38224 -1010 38229 -984
rect -18268 -1013 38229 -1010
rect 7089 -1031 7139 -1028
rect 7089 -1095 7092 -1031
rect 7136 -1095 7139 -1031
rect -17943 -1100 -17817 -1095
rect -17943 -1220 -17940 -1100
rect -17820 -1220 -17817 -1100
rect -17943 -1225 -17817 -1220
rect -15943 -1100 -15817 -1095
rect -15943 -1220 -15940 -1100
rect -15820 -1220 -15817 -1100
rect -15943 -1225 -15817 -1220
rect -13943 -1100 -13817 -1095
rect -13943 -1220 -13940 -1100
rect -13820 -1220 -13817 -1100
rect -13943 -1225 -13817 -1220
rect -11943 -1100 -11817 -1095
rect -11943 -1220 -11940 -1100
rect -11820 -1220 -11817 -1100
rect -11943 -1225 -11817 -1220
rect -9943 -1100 -9817 -1095
rect -9943 -1220 -9940 -1100
rect -9820 -1220 -9817 -1100
rect -9943 -1225 -9817 -1220
rect -7943 -1100 -7817 -1095
rect -7943 -1220 -7940 -1100
rect -7820 -1220 -7817 -1100
rect -7943 -1225 -7817 -1220
rect -5943 -1100 -5817 -1095
rect -5943 -1220 -5940 -1100
rect -5820 -1220 -5817 -1100
rect -5943 -1225 -5817 -1220
rect -3943 -1100 -3817 -1095
rect -3943 -1220 -3940 -1100
rect -3820 -1220 -3817 -1100
rect -3943 -1225 -3817 -1220
rect -1943 -1100 -1817 -1095
rect -1943 -1220 -1940 -1100
rect -1820 -1220 -1817 -1100
rect -1943 -1225 -1817 -1220
rect 57 -1100 183 -1095
rect 57 -1220 60 -1100
rect 180 -1220 183 -1100
rect 57 -1225 183 -1220
rect 1352 -1100 1478 -1095
rect 1352 -1220 1355 -1100
rect 1475 -1220 1478 -1100
rect 1352 -1225 1478 -1220
rect 6352 -1100 6478 -1095
rect 6352 -1220 6355 -1100
rect 6475 -1220 6478 -1100
rect 6352 -1225 6478 -1220
rect 7089 -1100 7478 -1095
rect 7089 -1220 7355 -1100
rect 7475 -1220 7478 -1100
rect 7089 -1225 7478 -1220
rect 19773 -1100 19899 -1095
rect 19773 -1220 19776 -1100
rect 19896 -1220 19899 -1100
rect 19773 -1225 19899 -1220
rect 21773 -1100 21899 -1095
rect 21773 -1220 21776 -1100
rect 21896 -1220 21899 -1100
rect 21773 -1225 21899 -1220
rect 23773 -1100 23899 -1095
rect 23773 -1220 23776 -1100
rect 23896 -1220 23899 -1100
rect 23773 -1225 23899 -1220
rect 25773 -1100 25899 -1095
rect 25773 -1220 25776 -1100
rect 25896 -1220 25899 -1100
rect 25773 -1225 25899 -1220
rect 27773 -1100 27899 -1095
rect 27773 -1220 27776 -1100
rect 27896 -1220 27899 -1100
rect 27773 -1225 27899 -1220
rect 29773 -1100 29899 -1095
rect 29773 -1220 29776 -1100
rect 29896 -1220 29899 -1100
rect 29773 -1225 29899 -1220
rect 31773 -1100 31899 -1095
rect 31773 -1220 31776 -1100
rect 31896 -1220 31899 -1100
rect 31773 -1225 31899 -1220
rect 33773 -1100 33899 -1095
rect 33773 -1220 33776 -1100
rect 33896 -1220 33899 -1100
rect 33773 -1225 33899 -1220
rect 35773 -1100 35899 -1095
rect 35773 -1220 35776 -1100
rect 35896 -1220 35899 -1100
rect 35773 -1225 35899 -1220
rect 37773 -1100 37899 -1095
rect 37773 -1220 37776 -1100
rect 37896 -1220 37899 -1100
rect 37773 -1225 37899 -1220
rect -18443 -1710 -18313 -1705
rect -18443 -1830 -18438 -1710
rect -18318 -1830 -18313 -1710
rect -18443 -1835 -18313 -1830
rect -16443 -1710 -16313 -1705
rect -16443 -1830 -16438 -1710
rect -16318 -1830 -16313 -1710
rect -16443 -1835 -16313 -1830
rect -14443 -1710 -14313 -1705
rect -14443 -1830 -14438 -1710
rect -14318 -1830 -14313 -1710
rect -14443 -1835 -14313 -1830
rect -12443 -1710 -12313 -1705
rect -12443 -1830 -12438 -1710
rect -12318 -1830 -12313 -1710
rect -12443 -1835 -12313 -1830
rect -10443 -1710 -10313 -1705
rect -10443 -1830 -10438 -1710
rect -10318 -1830 -10313 -1710
rect -10443 -1835 -10313 -1830
rect -8443 -1710 -8313 -1705
rect -8443 -1830 -8438 -1710
rect -8318 -1830 -8313 -1710
rect -8443 -1835 -8313 -1830
rect -6443 -1710 -6313 -1705
rect -6443 -1830 -6438 -1710
rect -6318 -1830 -6313 -1710
rect -6443 -1835 -6313 -1830
rect -4443 -1710 -4313 -1705
rect -4443 -1830 -4438 -1710
rect -4318 -1830 -4313 -1710
rect -4443 -1835 -4313 -1830
rect -2443 -1710 -2313 -1705
rect -2443 -1830 -2438 -1710
rect -2318 -1830 -2313 -1710
rect -2443 -1835 -2313 -1830
rect -443 -1710 -313 -1705
rect -443 -1830 -438 -1710
rect -318 -1830 -313 -1710
rect -443 -1835 -313 -1830
rect 852 -1710 982 -1705
rect 852 -1830 857 -1710
rect 977 -1830 982 -1710
rect 852 -1835 982 -1830
rect 5852 -1710 5982 -1705
rect 5852 -1830 5857 -1710
rect 5977 -1830 5982 -1710
rect 5852 -1835 5982 -1830
rect 6852 -1710 6982 -1705
rect 6852 -1830 6857 -1710
rect 6977 -1830 6982 -1710
rect 6852 -1835 6982 -1830
rect 20255 -1710 20385 -1705
rect 20255 -1830 20260 -1710
rect 20380 -1830 20385 -1710
rect 20255 -1835 20385 -1830
rect 22255 -1710 22385 -1705
rect 22255 -1830 22260 -1710
rect 22380 -1830 22385 -1710
rect 22255 -1835 22385 -1830
rect 24255 -1710 24385 -1705
rect 24255 -1830 24260 -1710
rect 24380 -1830 24385 -1710
rect 24255 -1835 24385 -1830
rect 26255 -1710 26385 -1705
rect 26255 -1830 26260 -1710
rect 26380 -1830 26385 -1710
rect 26255 -1835 26385 -1830
rect 28255 -1710 28385 -1705
rect 28255 -1830 28260 -1710
rect 28380 -1830 28385 -1710
rect 28255 -1835 28385 -1830
rect 30255 -1710 30385 -1705
rect 30255 -1830 30260 -1710
rect 30380 -1830 30385 -1710
rect 30255 -1835 30385 -1830
rect 32255 -1710 32385 -1705
rect 32255 -1830 32260 -1710
rect 32380 -1830 32385 -1710
rect 32255 -1835 32385 -1830
rect 34255 -1710 34385 -1705
rect 34255 -1830 34260 -1710
rect 34380 -1830 34385 -1710
rect 34255 -1835 34385 -1830
rect 36255 -1710 36385 -1705
rect 36255 -1830 36260 -1710
rect 36380 -1830 36385 -1710
rect 36255 -1835 36385 -1830
rect 38255 -1710 38385 -1705
rect 38255 -1830 38260 -1710
rect 38380 -1830 38385 -1710
rect 38255 -1835 38385 -1830
rect 4400 -2010 4800 -2000
rect 4400 -2190 4410 -2010
rect 4790 -2190 4800 -2010
rect 4400 -2200 4800 -2190
rect 17200 -2020 17800 -2000
rect 17200 -2180 17220 -2020
rect 17780 -2180 17800 -2020
rect 17200 -2200 17800 -2180
<< via2 >>
rect 2863 44215 3055 44259
rect 43 43733 435 43817
rect 19523 43733 19915 43817
rect 10923 42777 11113 42867
rect 2863 42715 3055 42759
rect 10655 42639 10845 42729
rect 10387 42501 10577 42591
rect 10119 42363 10309 42453
rect 43 42233 435 42317
rect 9851 42225 10041 42315
rect 19523 42233 19915 42317
rect 5325 41957 5815 42047
rect 14145 41957 14635 42047
rect 5325 41787 5815 41877
rect 14145 41787 14635 41877
rect 2863 41215 3055 41259
rect 43 40733 435 40817
rect 19523 40733 19915 40817
rect 2863 39715 3055 39759
rect 43 39233 435 39317
rect 19523 39233 19915 39317
rect 2863 38215 3055 38259
rect 43 37733 435 37817
rect 19523 37733 19915 37817
rect 2863 36915 3055 36959
rect 43 36233 435 36317
rect 19523 36233 19915 36317
rect 2863 35315 3055 35359
rect 43 34733 435 34817
rect 19523 34733 19915 34817
rect 2863 33715 3055 33759
rect 43 33233 435 33317
rect 19523 33233 19915 33317
rect 2863 32215 3055 32259
rect 43 31733 435 31817
rect 19523 31733 19915 31817
rect 2863 30915 3055 30959
rect 43 30233 435 30317
rect 19523 30233 19915 30317
rect 2863 29215 3055 29259
rect 3853 29447 4257 29451
rect 3853 29073 4257 29447
rect 3853 29047 4257 29073
rect 15703 29447 16107 29451
rect 15703 29073 16107 29447
rect 15703 29047 16107 29073
rect 5175 28997 5815 28998
rect 5175 28908 5815 28997
rect 14145 28997 14785 28998
rect 14145 28908 14785 28997
rect 43 28733 435 28817
rect 19523 28733 19915 28817
rect 2863 27715 3055 27759
rect 43 27233 435 27317
rect 19523 27233 19915 27317
rect 2863 26215 3055 26259
rect 43 25733 435 25817
rect 19523 25733 19915 25817
rect 2863 24715 3055 24759
rect 43 24233 435 24317
rect 19523 24233 19915 24317
rect 2863 23215 3055 23259
rect 43 22733 435 22817
rect 19523 22733 19915 22817
rect 2863 21715 3055 21759
rect 43 21233 435 21317
rect 5175 21105 5815 21295
rect 14145 21105 14785 21295
rect 19523 21233 19915 21317
rect 2863 20215 3055 20259
rect 43 19563 435 19817
rect 19523 19563 19915 19817
rect 10970 19340 11090 19460
rect 2863 18715 3055 18759
rect 43 18233 435 18317
rect 11070 18250 11190 18370
rect 19523 18233 19915 18317
rect 2863 17215 3055 17259
rect 43 16733 435 16817
rect 19523 16733 19915 16817
rect 2863 15715 3055 15759
rect 43 15233 435 15317
rect 19523 15233 19915 15317
rect 2863 14215 3055 14259
rect 43 13733 435 13817
rect 19523 13733 19915 13817
rect 2863 12715 3055 12759
rect 43 12233 435 12317
rect 19523 12233 19915 12317
rect 2863 11215 3055 11259
rect 43 10733 435 10817
rect 19523 10733 19915 10817
rect 2863 9715 3055 9759
rect 43 9233 435 9317
rect 19523 9233 19915 9317
rect 2863 8215 3055 8259
rect 43 7733 435 7817
rect 19523 7733 19915 7817
rect 2863 6715 3055 6759
rect 43 6233 435 6317
rect 19523 6233 19915 6317
rect 8779 6109 8969 6199
rect 9047 5941 9237 6031
rect 9315 5773 9505 5863
rect 9583 5605 9773 5695
rect 2863 5215 3055 5259
rect 43 4733 435 4817
rect 19523 4733 19915 4817
rect 2863 3715 3055 3759
rect 43 3233 435 3317
rect 19523 3233 19915 3317
rect 2863 2215 3055 2259
rect 43 1733 435 1817
rect 14903 2135 15097 2625
rect 14143 1585 14337 2075
rect 19523 1733 19915 1817
rect 2863 715 3055 759
rect 15675 595 16325 985
rect 40100 712 40220 832
rect 43 233 435 317
rect 19523 233 19915 317
rect -18215 -75 -18145 -5
rect -16215 -75 -16145 -5
rect -14215 -75 -14145 -5
rect -12215 -75 -12145 -5
rect -10215 -75 -10145 -5
rect -8215 -75 -8145 -5
rect -6215 -75 -6145 -5
rect -4215 -75 -4145 -5
rect -2215 -75 -2145 -5
rect -215 -75 -145 -5
rect 20105 -75 20175 -5
rect 22105 -75 22175 -5
rect 24105 -75 24175 -5
rect 26105 -75 26175 -5
rect 28105 -75 28175 -5
rect 30105 -75 30175 -5
rect 32105 -75 32175 -5
rect 34105 -75 34175 -5
rect 36105 -75 36175 -5
rect 38105 -75 38175 -5
rect -17940 -1220 -17820 -1100
rect -15940 -1220 -15820 -1100
rect -13940 -1220 -13820 -1100
rect -11940 -1220 -11820 -1100
rect -9940 -1220 -9820 -1100
rect -7940 -1220 -7820 -1100
rect -5940 -1220 -5820 -1100
rect -3940 -1220 -3820 -1100
rect -1940 -1220 -1820 -1100
rect 60 -1220 180 -1100
rect 1355 -1220 1475 -1100
rect 6355 -1220 6475 -1100
rect 7355 -1220 7475 -1100
rect 19776 -1220 19896 -1100
rect 21776 -1220 21896 -1100
rect 23776 -1220 23896 -1100
rect 25776 -1220 25896 -1100
rect 27776 -1220 27896 -1100
rect 29776 -1220 29896 -1100
rect 31776 -1220 31896 -1100
rect 33776 -1220 33896 -1100
rect 35776 -1220 35896 -1100
rect 37776 -1220 37896 -1100
rect -18438 -1830 -18318 -1710
rect -16438 -1830 -16318 -1710
rect -14438 -1830 -14318 -1710
rect -12438 -1830 -12318 -1710
rect -10438 -1830 -10318 -1710
rect -8438 -1830 -8318 -1710
rect -6438 -1830 -6318 -1710
rect -4438 -1830 -4318 -1710
rect -2438 -1830 -2318 -1710
rect -438 -1830 -318 -1710
rect 857 -1830 977 -1710
rect 5857 -1830 5977 -1710
rect 6857 -1830 6977 -1710
rect 20260 -1830 20380 -1710
rect 22260 -1830 22380 -1710
rect 24260 -1830 24380 -1710
rect 26260 -1830 26380 -1710
rect 28260 -1830 28380 -1710
rect 30260 -1830 30380 -1710
rect 32260 -1830 32380 -1710
rect 34260 -1830 34380 -1710
rect 36260 -1830 36380 -1710
rect 38260 -1830 38380 -1710
rect 4410 -2190 4790 -2010
rect 17220 -2180 17780 -2020
<< metal3 >>
rect 2860 44259 3520 44605
rect 2860 44215 2863 44259
rect 3055 44215 3520 44259
rect 40 43817 440 43820
rect 40 43733 43 43817
rect 435 43733 440 43817
rect 40 42317 440 43733
rect 40 42233 43 42317
rect 435 42233 440 42317
rect 40 40817 440 42233
rect 40 40733 43 40817
rect 435 40733 440 40817
rect 40 39317 440 40733
rect 40 39233 43 39317
rect 435 39233 440 39317
rect 40 37817 440 39233
rect 40 37733 43 37817
rect 435 37733 440 37817
rect 40 36317 440 37733
rect 40 36233 43 36317
rect 435 36233 440 36317
rect 40 34817 440 36233
rect 40 34733 43 34817
rect 435 34733 440 34817
rect 40 33317 440 34733
rect 40 33233 43 33317
rect 435 33233 440 33317
rect 40 31817 440 33233
rect 40 31733 43 31817
rect 435 31733 440 31817
rect 40 30317 440 31733
rect 40 30233 43 30317
rect 435 30233 440 30317
rect 40 28817 440 30233
rect 40 28733 43 28817
rect 435 28733 440 28817
rect 40 27317 440 28733
rect 40 27233 43 27317
rect 435 27233 440 27317
rect 40 25817 440 27233
rect 40 25733 43 25817
rect 435 25733 440 25817
rect 40 24317 440 25733
rect 40 24233 43 24317
rect 435 24233 440 24317
rect 40 22817 440 24233
rect 40 22733 43 22817
rect 435 22733 440 22817
rect 40 21317 440 22733
rect 40 21233 43 21317
rect 435 21233 440 21317
rect 40 19817 440 21233
rect 40 19563 43 19817
rect 435 19563 440 19817
rect 40 18317 440 19563
rect 40 18233 43 18317
rect 435 18233 440 18317
rect 40 16817 440 18233
rect 40 16733 43 16817
rect 435 16733 440 16817
rect 40 15317 440 16733
rect 40 15233 43 15317
rect 435 15233 440 15317
rect 40 13817 440 15233
rect 40 13733 43 13817
rect 435 13733 440 13817
rect 40 12317 440 13733
rect 40 12233 43 12317
rect 435 12233 440 12317
rect 40 10817 440 12233
rect 40 10733 43 10817
rect 435 10733 440 10817
rect 40 9317 440 10733
rect 40 9233 43 9317
rect 435 9233 440 9317
rect 40 7817 440 9233
rect 40 7733 43 7817
rect 435 7733 440 7817
rect 40 6317 440 7733
rect 40 6233 43 6317
rect 435 6233 440 6317
rect 40 4817 440 6233
rect 40 4733 43 4817
rect 435 4733 440 4817
rect 40 3317 440 4733
rect 40 3233 43 3317
rect 435 3233 440 3317
rect 40 1817 440 3233
rect 40 1733 43 1817
rect 435 1733 440 1817
rect 40 317 440 1733
rect 40 233 43 317
rect 435 233 440 317
rect 40 230 440 233
rect 2860 42759 3520 44215
rect 2860 42715 2863 42759
rect 3055 42715 3520 42759
rect 2860 41259 3520 42715
rect 4100 44300 4900 45600
rect 4100 43930 4130 44300
rect 4870 43930 4900 44300
rect 4100 42800 4900 43930
rect 6100 44800 6900 45600
rect 6100 44430 6130 44800
rect 6870 44430 6900 44800
rect 4100 42047 5900 42800
rect 4100 42000 5325 42047
rect 4400 41957 5325 42000
rect 5815 41957 5900 42047
rect 4400 41950 5900 41957
rect 2860 41215 2863 41259
rect 3055 41215 3520 41259
rect 2860 39759 3520 41215
rect 2860 39715 2863 39759
rect 3055 39715 3520 39759
rect 2860 38259 3520 39715
rect 2860 38215 2863 38259
rect 3055 38215 3520 38259
rect 2860 36959 3520 38215
rect 2860 36915 2863 36959
rect 3055 36915 3520 36959
rect 2860 35359 3520 36915
rect 2860 35315 2863 35359
rect 3055 35315 3520 35359
rect 2860 33759 3520 35315
rect 2860 33715 2863 33759
rect 3055 33715 3520 33759
rect 2860 32259 3520 33715
rect 2860 32215 2863 32259
rect 3055 32215 3520 32259
rect 2860 30959 3520 32215
rect 2860 30915 2863 30959
rect 3055 30915 3520 30959
rect 2860 29259 3520 30915
rect 2860 29215 2863 29259
rect 3055 29215 3520 29259
rect 2860 27759 3520 29215
rect 2860 27715 2863 27759
rect 3055 27715 3520 27759
rect 2860 26259 3520 27715
rect 2860 26215 2863 26259
rect 3055 26215 3520 26259
rect 2860 24759 3520 26215
rect 2860 24715 2863 24759
rect 3055 24715 3520 24759
rect 2860 23259 3520 24715
rect 2860 23215 2863 23259
rect 3055 23215 3520 23259
rect 2860 21759 3520 23215
rect 2860 21715 2863 21759
rect 3055 21715 3520 21759
rect 2860 20259 3520 21715
rect 2860 20215 2863 20259
rect 3055 20215 3520 20259
rect 2860 18759 3520 20215
rect 2860 18715 2863 18759
rect 3055 18715 3520 18759
rect 2860 17259 3520 18715
rect 2860 17215 2863 17259
rect 3055 17215 3520 17259
rect 2860 15759 3520 17215
rect 2860 15715 2863 15759
rect 3055 15715 3520 15759
rect 2860 14259 3520 15715
rect 2860 14215 2863 14259
rect 3055 14215 3520 14259
rect 2860 12759 3520 14215
rect 2860 12715 2863 12759
rect 3055 12715 3520 12759
rect 2860 11259 3520 12715
rect 2860 11215 2863 11259
rect 3055 11215 3520 11259
rect 2860 9759 3520 11215
rect 2860 9715 2863 9759
rect 3055 9715 3520 9759
rect 2860 8259 3520 9715
rect 2860 8215 2863 8259
rect 3055 8215 3520 8259
rect 2860 6759 3520 8215
rect 2860 6715 2863 6759
rect 3055 6715 3520 6759
rect 2860 5259 3520 6715
rect 2860 5215 2863 5259
rect 3055 5215 3520 5259
rect 2860 3759 3520 5215
rect 2860 3715 2863 3759
rect 3055 3715 3520 3759
rect 2860 2259 3520 3715
rect 2860 2215 2863 2259
rect 3055 2215 3520 2259
rect 2860 759 3520 2215
rect 2860 715 2863 759
rect 3055 715 3520 759
rect 100 80 800 100
rect -18600 -200 -18400 0
rect -18220 -5 -18140 0
rect -18220 -75 -18215 -5
rect -18145 -75 -18140 -5
rect -18220 -80 -18140 -75
rect -16600 -200 -16400 0
rect -16220 -5 -16140 0
rect -16220 -75 -16215 -5
rect -16145 -75 -16140 -5
rect -16220 -80 -16140 -75
rect -14600 -200 -14400 0
rect -14220 -5 -14140 0
rect -14220 -75 -14215 -5
rect -14145 -75 -14140 -5
rect -14220 -80 -14140 -75
rect -12600 -200 -12400 0
rect -12220 -5 -12140 0
rect -12220 -75 -12215 -5
rect -12145 -75 -12140 -5
rect -12220 -80 -12140 -75
rect -10600 -200 -10400 0
rect -10220 -5 -10140 0
rect -10220 -75 -10215 -5
rect -10145 -75 -10140 -5
rect -10220 -80 -10140 -75
rect -8600 -200 -8400 0
rect -8220 -5 -8140 0
rect -8220 -75 -8215 -5
rect -8145 -75 -8140 -5
rect -8220 -80 -8140 -75
rect -6600 -200 -6400 0
rect -6220 -5 -6140 0
rect -6220 -75 -6215 -5
rect -6145 -75 -6140 -5
rect -6220 -80 -6140 -75
rect -4600 -200 -4400 0
rect -4220 -5 -4140 0
rect -4220 -75 -4215 -5
rect -4145 -75 -4140 -5
rect -4220 -80 -4140 -75
rect -2600 -200 -2400 0
rect -2220 -5 -2140 0
rect -2220 -75 -2215 -5
rect -2145 -75 -2140 -5
rect -2220 -80 -2140 -75
rect -600 -200 -400 0
rect -220 -5 -140 0
rect -220 -75 -215 -5
rect -145 -75 -140 -5
rect -220 -80 -140 -75
rect 100 -200 120 80
rect -18600 -380 120 -200
rect 780 -380 800 80
rect -18600 -600 800 -380
rect 2090 80 2750 100
rect 2090 -380 2110 80
rect 2730 -380 2750 80
rect -17943 -1100 -17817 -1097
rect -17943 -1220 -17940 -1100
rect -17820 -1220 -17817 -1100
rect -17943 -1223 -17817 -1220
rect -15943 -1100 -15817 -1097
rect -15943 -1220 -15940 -1100
rect -15820 -1220 -15817 -1100
rect -15943 -1223 -15817 -1220
rect -13943 -1100 -13817 -1097
rect -13943 -1220 -13940 -1100
rect -13820 -1220 -13817 -1100
rect -13943 -1223 -13817 -1220
rect -11943 -1100 -11817 -1097
rect -11943 -1220 -11940 -1100
rect -11820 -1220 -11817 -1100
rect -11943 -1223 -11817 -1220
rect -9943 -1100 -9817 -1097
rect -9943 -1220 -9940 -1100
rect -9820 -1220 -9817 -1100
rect -9943 -1223 -9817 -1220
rect -7943 -1100 -7817 -1097
rect -7943 -1220 -7940 -1100
rect -7820 -1220 -7817 -1100
rect -7943 -1223 -7817 -1220
rect -5943 -1100 -5817 -1097
rect -5943 -1220 -5940 -1100
rect -5820 -1220 -5817 -1100
rect -5943 -1223 -5817 -1220
rect -3943 -1100 -3817 -1097
rect -3943 -1220 -3940 -1100
rect -3820 -1220 -3817 -1100
rect -3943 -1223 -3817 -1220
rect -1943 -1100 -1817 -1097
rect -1943 -1220 -1940 -1100
rect -1820 -1220 -1817 -1100
rect -1943 -1223 -1817 -1220
rect 57 -1100 183 -1097
rect 57 -1220 60 -1100
rect 180 -1220 183 -1100
rect 57 -1223 183 -1220
rect 1352 -1100 1478 -1097
rect 1352 -1220 1355 -1100
rect 1475 -1220 1478 -1100
rect 1352 -1223 1478 -1220
rect -18443 -1710 -18313 -1705
rect -18443 -1830 -18438 -1710
rect -18318 -1830 -18313 -1710
rect -18443 -1835 -18313 -1830
rect -16443 -1710 -16313 -1705
rect -16443 -1830 -16438 -1710
rect -16318 -1830 -16313 -1710
rect -16443 -1835 -16313 -1830
rect -14443 -1710 -14313 -1705
rect -14443 -1830 -14438 -1710
rect -14318 -1830 -14313 -1710
rect -14443 -1835 -14313 -1830
rect -12443 -1710 -12313 -1705
rect -12443 -1830 -12438 -1710
rect -12318 -1830 -12313 -1710
rect -12443 -1835 -12313 -1830
rect -10443 -1710 -10313 -1705
rect -10443 -1830 -10438 -1710
rect -10318 -1830 -10313 -1710
rect -10443 -1835 -10313 -1830
rect -8443 -1710 -8313 -1705
rect -8443 -1830 -8438 -1710
rect -8318 -1830 -8313 -1710
rect -8443 -1835 -8313 -1830
rect -6443 -1710 -6313 -1705
rect -6443 -1830 -6438 -1710
rect -6318 -1830 -6313 -1710
rect -6443 -1835 -6313 -1830
rect -4443 -1710 -4313 -1705
rect -4443 -1830 -4438 -1710
rect -4318 -1830 -4313 -1710
rect -4443 -1835 -4313 -1830
rect -2443 -1710 -2313 -1705
rect -2443 -1830 -2438 -1710
rect -2318 -1830 -2313 -1710
rect -2443 -1835 -2313 -1830
rect -443 -1710 -313 -1705
rect -443 -1830 -438 -1710
rect -318 -1830 -313 -1710
rect -443 -1835 -313 -1830
rect 852 -1710 982 -1705
rect 852 -1830 857 -1710
rect 977 -1830 982 -1710
rect 852 -1835 982 -1830
rect 2090 -2600 2750 -380
rect 2860 -2600 3520 715
rect 3630 29451 4290 41530
rect 3630 29047 3853 29451
rect 4257 29047 4290 29451
rect 3630 18397 4290 29047
rect 3630 17403 3633 18397
rect 4287 17403 4290 18397
rect 3630 -1703 4290 17403
rect 4400 700 5060 41950
rect 6100 41900 6900 44430
rect 7300 43600 7500 45600
rect 7900 43900 8100 45600
rect 8500 44200 8700 45600
rect 9100 44500 9300 45600
rect 9700 44800 9900 45600
rect 9700 44600 10046 44800
rect 10300 44620 10500 45600
rect 9100 44300 9778 44500
rect 8500 44000 9510 44200
rect 7900 43700 9242 43900
rect 7300 43400 8974 43600
rect 5170 41877 6900 41900
rect 5170 41787 5325 41877
rect 5815 41787 6900 41877
rect 5170 41100 6900 41787
rect 5170 28998 5820 41100
rect 5170 28908 5175 28998
rect 5815 28908 5820 28998
rect 5170 21295 5820 28908
rect 5170 21105 5175 21295
rect 5815 21105 5820 21295
rect 5170 20330 5200 21105
rect 5790 20330 5820 21105
rect 5170 -503 5820 20330
rect 8774 6199 8974 43400
rect 8774 6109 8779 6199
rect 8969 6109 8974 6199
rect 8774 6104 8974 6109
rect 9042 6031 9242 43700
rect 9042 5941 9047 6031
rect 9237 5941 9242 6031
rect 9042 5936 9242 5941
rect 9310 5863 9510 44000
rect 9310 5773 9315 5863
rect 9505 5773 9510 5863
rect 9310 5768 9510 5773
rect 9578 5695 9778 44300
rect 9846 42315 10046 44600
rect 10114 44420 10500 44620
rect 10114 42453 10314 44420
rect 10900 44320 11100 45600
rect 10382 44120 11100 44320
rect 10382 42591 10582 44120
rect 11500 44020 11700 45600
rect 10650 43820 11700 44020
rect 10650 42729 10850 43820
rect 12100 43720 12300 45600
rect 10918 43520 12300 43720
rect 12700 44300 13500 45600
rect 14700 44800 15500 45600
rect 14700 44430 14730 44800
rect 15470 44430 15500 44800
rect 14700 44420 15500 44430
rect 12700 43930 12730 44300
rect 13470 43930 13500 44300
rect 10918 42867 11118 43520
rect 10918 42777 10923 42867
rect 11113 42777 11118 42867
rect 10918 42772 11118 42777
rect 10650 42639 10655 42729
rect 10845 42639 10850 42729
rect 10650 42634 10850 42639
rect 12700 42750 13500 43930
rect 19520 43817 19920 43820
rect 19520 43733 19523 43817
rect 19915 43733 19920 43817
rect 10382 42501 10387 42591
rect 10577 42501 10582 42591
rect 10382 42496 10582 42501
rect 10114 42363 10119 42453
rect 10309 42363 10314 42453
rect 10114 42358 10314 42363
rect 9846 42225 9851 42315
rect 10041 42225 10046 42315
rect 9846 42220 10046 42225
rect 12700 42047 15560 42750
rect 12700 41957 14145 42047
rect 14635 41957 15560 42047
rect 12700 41950 15560 41957
rect 13700 41880 14800 41890
rect 13700 41710 13710 41880
rect 14490 41877 14800 41880
rect 14635 41787 14800 41877
rect 14490 41710 14800 41787
rect 13700 41700 14800 41710
rect 14140 41100 14800 41700
rect 14140 28998 14790 41100
rect 14140 28908 14145 28998
rect 14785 28908 14790 28998
rect 14140 21295 14790 28908
rect 14140 21105 14145 21295
rect 14785 21105 14790 21295
rect 10965 20427 11095 20430
rect 10965 20303 10968 20427
rect 11092 20303 11095 20427
rect 10965 19460 11095 20303
rect 10965 19340 10970 19460
rect 11090 19340 11095 19460
rect 10965 19335 11095 19340
rect 14140 20330 14170 21105
rect 14760 20330 14790 21105
rect 11065 18370 11195 18375
rect 11065 18250 11070 18370
rect 11190 18250 11195 18370
rect 11065 18245 11195 18250
rect 9578 5605 9583 5695
rect 9773 5605 9778 5695
rect 9578 5600 9778 5605
rect 5170 -1497 5173 -503
rect 5817 -1497 5820 -503
rect 14140 2075 14790 20330
rect 14140 1585 14143 2075
rect 14337 1585 14790 2075
rect 14140 -503 14790 1585
rect 14900 2625 15560 41950
rect 19520 42317 19920 43733
rect 19520 42233 19523 42317
rect 19915 42233 19920 42317
rect 14900 2135 14903 2625
rect 15097 2135 15560 2625
rect 14900 1077 15560 2135
rect 15670 29451 16330 41570
rect 15670 29047 15703 29451
rect 16107 29047 16330 29451
rect 15670 18397 16330 29047
rect 15670 17403 15673 18397
rect 16327 17403 16330 18397
rect 6352 -1100 6478 -1097
rect 6352 -1220 6355 -1100
rect 6475 -1220 6478 -1100
rect 6352 -1223 6478 -1220
rect 7352 -1100 7478 -1097
rect 7352 -1220 7355 -1100
rect 7475 -1220 7478 -1100
rect 7352 -1223 7478 -1220
rect 5170 -1500 5820 -1497
rect 14140 -1497 14143 -503
rect 14787 -1497 14790 -503
rect 14140 -1500 14790 -1497
rect 15670 985 16330 17403
rect 15670 595 15675 985
rect 16325 595 16330 985
rect 3630 -2297 3633 -1703
rect 4287 -2297 4290 -1703
rect 15670 -1703 16330 595
rect 19520 40817 19920 42233
rect 19520 40733 19523 40817
rect 19915 40733 19920 40817
rect 19520 39317 19920 40733
rect 19520 39233 19523 39317
rect 19915 39233 19920 39317
rect 19520 37817 19920 39233
rect 19520 37733 19523 37817
rect 19915 37733 19920 37817
rect 19520 36317 19920 37733
rect 19520 36233 19523 36317
rect 19915 36233 19920 36317
rect 19520 34817 19920 36233
rect 19520 34733 19523 34817
rect 19915 34733 19920 34817
rect 19520 33317 19920 34733
rect 19520 33233 19523 33317
rect 19915 33233 19920 33317
rect 19520 31817 19920 33233
rect 19520 31733 19523 31817
rect 19915 31733 19920 31817
rect 19520 30317 19920 31733
rect 19520 30233 19523 30317
rect 19915 30233 19920 30317
rect 19520 28817 19920 30233
rect 19520 28733 19523 28817
rect 19915 28733 19920 28817
rect 19520 27317 19920 28733
rect 19520 27233 19523 27317
rect 19915 27233 19920 27317
rect 19520 25817 19920 27233
rect 19520 25733 19523 25817
rect 19915 25733 19920 25817
rect 19520 24317 19920 25733
rect 19520 24233 19523 24317
rect 19915 24233 19920 24317
rect 19520 22817 19920 24233
rect 19520 22733 19523 22817
rect 19915 22733 19920 22817
rect 19520 21317 19920 22733
rect 19520 21233 19523 21317
rect 19915 21233 19920 21317
rect 19520 19817 19920 21233
rect 19520 19563 19523 19817
rect 19915 19563 19920 19817
rect 19520 18317 19920 19563
rect 19520 18233 19523 18317
rect 19915 18233 19920 18317
rect 19520 16817 19920 18233
rect 19520 16733 19523 16817
rect 19915 16733 19920 16817
rect 19520 15317 19920 16733
rect 19520 15233 19523 15317
rect 19915 15233 19920 15317
rect 19520 13817 19920 15233
rect 19520 13733 19523 13817
rect 19915 13733 19920 13817
rect 19520 12317 19920 13733
rect 19520 12233 19523 12317
rect 19915 12233 19920 12317
rect 19520 10817 19920 12233
rect 19520 10733 19523 10817
rect 19915 10733 19920 10817
rect 19520 9317 19920 10733
rect 19520 9233 19523 9317
rect 19915 9233 19920 9317
rect 19520 7817 19920 9233
rect 19520 7733 19523 7817
rect 19915 7733 19920 7817
rect 19520 6317 19920 7733
rect 19520 6233 19523 6317
rect 19915 6233 19920 6317
rect 19520 4817 19920 6233
rect 19520 4733 19523 4817
rect 19915 4733 19920 4817
rect 19520 3317 19920 4733
rect 19520 3233 19523 3317
rect 19915 3233 19920 3317
rect 19520 1817 19920 3233
rect 19520 1733 19523 1817
rect 19915 1733 19920 1817
rect 19520 317 19920 1733
rect 40093 832 40242 849
rect 40093 712 40100 832
rect 40220 712 40242 832
rect 40093 705 40242 712
rect 19520 233 19523 317
rect 19915 233 19920 317
rect 19520 230 19920 233
rect 19160 70 19860 100
rect 19160 -370 19190 70
rect 19830 -200 19860 70
rect 20100 -5 20180 0
rect 20100 -75 20105 -5
rect 20175 -75 20180 -5
rect 20100 -80 20180 -75
rect 20360 -200 20560 0
rect 22100 -5 22180 0
rect 22100 -75 22105 -5
rect 22175 -75 22180 -5
rect 22100 -80 22180 -75
rect 22360 -200 22560 0
rect 24100 -5 24180 0
rect 24100 -75 24105 -5
rect 24175 -75 24180 -5
rect 24100 -80 24180 -75
rect 24360 -200 24560 0
rect 26100 -5 26180 0
rect 26100 -75 26105 -5
rect 26175 -75 26180 -5
rect 26100 -80 26180 -75
rect 26360 -200 26560 0
rect 28100 -5 28180 0
rect 28100 -75 28105 -5
rect 28175 -75 28180 -5
rect 28100 -80 28180 -75
rect 28360 -200 28560 0
rect 30100 -5 30180 0
rect 30100 -75 30105 -5
rect 30175 -75 30180 -5
rect 30100 -80 30180 -75
rect 30360 -200 30560 0
rect 32100 -5 32180 0
rect 32100 -75 32105 -5
rect 32175 -75 32180 -5
rect 32100 -80 32180 -75
rect 32360 -200 32560 0
rect 34100 -5 34180 0
rect 34100 -75 34105 -5
rect 34175 -75 34180 -5
rect 34100 -80 34180 -75
rect 34360 -200 34560 0
rect 36100 -5 36180 0
rect 36100 -75 36105 -5
rect 36175 -75 36180 -5
rect 36100 -80 36180 -75
rect 36360 -200 36560 0
rect 38100 -5 38180 0
rect 38100 -75 38105 -5
rect 38175 -75 38180 -5
rect 38100 -80 38180 -75
rect 38360 -200 38560 0
rect 19830 -370 38560 -200
rect 19160 -600 38560 -370
rect 24500 -720 26100 -700
rect 19773 -1100 19899 -1097
rect 19773 -1220 19776 -1100
rect 19896 -1220 19899 -1100
rect 19773 -1223 19899 -1220
rect 21773 -1100 21899 -1097
rect 21773 -1220 21776 -1100
rect 21896 -1220 21899 -1100
rect 21773 -1223 21899 -1220
rect 23773 -1100 23899 -1097
rect 23773 -1220 23776 -1100
rect 23896 -1220 23899 -1100
rect 23773 -1223 23899 -1220
rect 5852 -1710 5982 -1705
rect 5852 -1830 5857 -1710
rect 5977 -1830 5982 -1710
rect 5852 -1835 5982 -1830
rect 6852 -1710 6982 -1705
rect 6852 -1830 6857 -1710
rect 6977 -1830 6982 -1710
rect 6852 -1835 6982 -1830
rect 3630 -2300 4290 -2297
rect 4400 -2010 4800 -2000
rect 4400 -2190 4410 -2010
rect 4790 -2190 4800 -2010
rect 4400 -2600 4800 -2190
rect 15670 -2297 15673 -1703
rect 16327 -2297 16330 -1703
rect 24500 -1480 24520 -720
rect 26080 -1480 26100 -720
rect 27773 -1100 27899 -1097
rect 27773 -1220 27776 -1100
rect 27896 -1220 27899 -1100
rect 27773 -1223 27899 -1220
rect 29773 -1100 29899 -1097
rect 29773 -1220 29776 -1100
rect 29896 -1220 29899 -1100
rect 29773 -1223 29899 -1220
rect 31773 -1100 31899 -1097
rect 31773 -1220 31776 -1100
rect 31896 -1220 31899 -1100
rect 31773 -1223 31899 -1220
rect 33773 -1100 33899 -1097
rect 33773 -1220 33776 -1100
rect 33896 -1220 33899 -1100
rect 33773 -1223 33899 -1220
rect 35773 -1100 35899 -1097
rect 35773 -1220 35776 -1100
rect 35896 -1220 35899 -1100
rect 35773 -1223 35899 -1220
rect 37773 -1100 37899 -1097
rect 37773 -1220 37776 -1100
rect 37896 -1220 37899 -1100
rect 37773 -1223 37899 -1220
rect 20255 -1710 20385 -1705
rect 20255 -1830 20260 -1710
rect 20380 -1830 20385 -1710
rect 20255 -1835 20385 -1830
rect 22255 -1710 22385 -1705
rect 22255 -1830 22260 -1710
rect 22380 -1830 22385 -1710
rect 22255 -1835 22385 -1830
rect 24255 -1710 24385 -1705
rect 24255 -1830 24260 -1710
rect 24380 -1830 24385 -1710
rect 24255 -1835 24385 -1830
rect 15670 -2300 16330 -2297
rect 17190 -2020 17800 -2000
rect 17190 -2180 17220 -2020
rect 17780 -2180 17800 -2020
rect 17190 -2600 17800 -2180
rect 24500 -2400 26100 -1480
rect 26255 -1710 26385 -1705
rect 26255 -1830 26260 -1710
rect 26380 -1830 26385 -1710
rect 26255 -1835 26385 -1830
rect 28255 -1710 28385 -1705
rect 28255 -1830 28260 -1710
rect 28380 -1830 28385 -1710
rect 28255 -1835 28385 -1830
rect 30255 -1710 30385 -1705
rect 30255 -1830 30260 -1710
rect 30380 -1830 30385 -1710
rect 30255 -1835 30385 -1830
rect 32255 -1710 32385 -1705
rect 32255 -1830 32260 -1710
rect 32380 -1830 32385 -1710
rect 32255 -1835 32385 -1830
rect 34255 -1710 34385 -1705
rect 34255 -1830 34260 -1710
rect 34380 -1830 34385 -1710
rect 34255 -1835 34385 -1830
rect 36255 -1710 36385 -1705
rect 36255 -1830 36260 -1710
rect 36380 -1830 36385 -1710
rect 36255 -1835 36385 -1830
rect 38255 -1710 38385 -1705
rect 38255 -1830 38260 -1710
rect 38380 -1830 38385 -1710
rect 38255 -1835 38385 -1830
rect 23900 -2600 26100 -2400
<< via3 >>
rect 4130 43930 4870 44300
rect 6130 44430 6870 44800
rect 120 -380 780 80
rect 2110 -380 2730 80
rect -17940 -1220 -17820 -1100
rect -15940 -1220 -15820 -1100
rect -13940 -1220 -13820 -1100
rect -11940 -1220 -11820 -1100
rect -9940 -1220 -9820 -1100
rect -7940 -1220 -7820 -1100
rect -5940 -1220 -5820 -1100
rect -3940 -1220 -3820 -1100
rect -1940 -1220 -1820 -1100
rect 60 -1220 180 -1100
rect 1355 -1220 1475 -1100
rect -18438 -1830 -18318 -1710
rect -16438 -1830 -16318 -1710
rect -14438 -1830 -14318 -1710
rect -12438 -1830 -12318 -1710
rect -10438 -1830 -10318 -1710
rect -8438 -1830 -8318 -1710
rect -6438 -1830 -6318 -1710
rect -4438 -1830 -4318 -1710
rect -2438 -1830 -2318 -1710
rect -438 -1830 -318 -1710
rect 857 -1830 977 -1710
rect 3633 17403 4287 18397
rect 5200 21105 5790 21270
rect 5200 20330 5790 21105
rect 14730 44430 15470 44800
rect 12730 43930 13470 44300
rect 13710 41877 14490 41880
rect 13710 41787 14145 41877
rect 14145 41787 14490 41877
rect 13710 41710 14490 41787
rect 14170 21105 14760 21270
rect 10968 20303 11092 20427
rect 14170 20330 14760 21105
rect 11070 18250 11190 18370
rect 5173 -1497 5817 -503
rect 15673 17403 16327 18397
rect 6355 -1220 6475 -1100
rect 7355 -1220 7475 -1100
rect 14143 -1497 14787 -503
rect 3633 -2297 4287 -1703
rect 40100 712 40220 832
rect 19190 -370 19830 70
rect 19776 -1220 19896 -1100
rect 21776 -1220 21896 -1100
rect 23776 -1220 23896 -1100
rect 5857 -1830 5977 -1710
rect 6857 -1830 6977 -1710
rect 15673 -2297 16327 -1703
rect 24520 -1100 26080 -720
rect 24520 -1220 25776 -1100
rect 25776 -1220 25896 -1100
rect 25896 -1220 26080 -1100
rect 24520 -1480 26080 -1220
rect 27776 -1220 27896 -1100
rect 29776 -1220 29896 -1100
rect 31776 -1220 31896 -1100
rect 33776 -1220 33896 -1100
rect 35776 -1220 35896 -1100
rect 37776 -1220 37896 -1100
rect 20260 -1830 20380 -1710
rect 22260 -1830 22380 -1710
rect 24260 -1830 24380 -1710
rect 26260 -1830 26380 -1710
rect 28260 -1830 28380 -1710
rect 30260 -1830 30380 -1710
rect 32260 -1830 32380 -1710
rect 34260 -1830 34380 -1710
rect 36260 -1830 36380 -1710
rect 38260 -1830 38380 -1710
<< metal4 >>
rect 6100 44800 15500 44801
rect 6100 44430 6130 44800
rect 6870 44430 14730 44800
rect 15470 44430 15500 44800
rect 6100 44400 15500 44430
rect 4100 44300 4900 44301
rect 12700 44300 13500 44301
rect 40 18400 540 44300
rect 4100 43930 4130 44300
rect 4870 43930 12730 44300
rect 13470 43930 13500 44300
rect 4100 43900 13500 43930
rect 13700 41880 14500 44400
rect 13700 41710 13710 41880
rect 14490 41710 14500 41880
rect 13700 41700 14500 41710
rect 5170 21270 14790 21300
rect 5170 20330 5200 21270
rect 5790 20427 14170 21270
rect 5790 20330 10968 20427
rect 5170 20303 10968 20330
rect 11092 20330 14170 20427
rect 14760 20330 14790 21270
rect 11092 20303 14790 20330
rect 5170 20300 14790 20303
rect 19420 18400 19920 44300
rect 40 18397 19920 18400
rect 40 17403 3633 18397
rect 4287 18370 15673 18397
rect 4287 18250 11070 18370
rect 11190 18250 15673 18370
rect 4287 17403 15673 18250
rect 16327 17403 19920 18397
rect 40 17400 19920 17403
rect 40 400 540 17400
rect 19420 400 19920 17400
rect 40093 832 40242 849
rect 40093 712 40100 832
rect 40220 712 40242 832
rect 40093 705 40242 712
rect 100 80 19860 100
rect -18900 -500 -18300 -380
rect -16900 -500 -16300 -380
rect -14900 -500 -14300 -380
rect -12900 -500 -12300 -380
rect -10900 -500 -10300 -380
rect -8900 -500 -8300 -380
rect -6900 -500 -6300 -380
rect -4900 -500 -4300 -380
rect -2900 -500 -2300 -380
rect -900 -500 -300 -380
rect 100 -380 120 80
rect 780 -380 2110 80
rect 2730 70 19860 80
rect 2730 -370 19190 70
rect 19830 -370 19860 70
rect 2730 -380 19860 -370
rect 100 -400 19860 -380
rect 20260 -500 20860 -380
rect 22260 -500 22860 -380
rect 24260 -500 24860 -380
rect 26260 -500 26860 -380
rect 28260 -500 28860 -380
rect 30260 -500 30860 -380
rect 32260 -500 32860 -380
rect 34260 -500 34860 -380
rect 36260 -500 36860 -380
rect 38260 -500 38860 -380
rect -20500 -503 40460 -500
rect -20500 -520 5173 -503
rect -20500 -1480 -20480 -520
rect -20120 -1100 5173 -520
rect -20120 -1220 -17940 -1100
rect -17820 -1220 -15940 -1100
rect -15820 -1220 -13940 -1100
rect -13820 -1220 -11940 -1100
rect -11820 -1220 -9940 -1100
rect -9820 -1220 -7940 -1100
rect -7820 -1220 -5940 -1100
rect -5820 -1220 -3940 -1100
rect -3820 -1220 -1940 -1100
rect -1820 -1220 60 -1100
rect 180 -1220 1355 -1100
rect 1475 -1220 5173 -1100
rect -20120 -1480 5173 -1220
rect -20500 -1497 5173 -1480
rect 5817 -1100 14143 -503
rect 5817 -1220 6355 -1100
rect 6475 -1220 7355 -1100
rect 7475 -1220 14143 -1100
rect 5817 -1497 14143 -1220
rect 14787 -520 40460 -503
rect 14787 -720 40080 -520
rect 14787 -1100 24520 -720
rect 14787 -1220 19776 -1100
rect 19896 -1220 21776 -1100
rect 21896 -1220 23776 -1100
rect 23896 -1220 24520 -1100
rect 14787 -1480 24520 -1220
rect 26080 -1100 40080 -720
rect 26080 -1220 27776 -1100
rect 27896 -1220 29776 -1100
rect 29896 -1220 31776 -1100
rect 31896 -1220 33776 -1100
rect 33896 -1220 35776 -1100
rect 35896 -1220 37776 -1100
rect 37896 -1220 40080 -1100
rect 26080 -1480 40080 -1220
rect 40440 -1480 40460 -520
rect 14787 -1497 40460 -1480
rect -20500 -1500 40460 -1497
rect -18500 -1703 38390 -1700
rect -18500 -1710 3633 -1703
rect -18500 -1830 -18438 -1710
rect -18318 -1830 -16438 -1710
rect -16318 -1830 -14438 -1710
rect -14318 -1830 -12438 -1710
rect -12318 -1830 -10438 -1710
rect -10318 -1830 -8438 -1710
rect -8318 -1830 -6438 -1710
rect -6318 -1830 -4438 -1710
rect -4318 -1830 -2438 -1710
rect -2318 -1830 -438 -1710
rect -318 -1830 857 -1710
rect 977 -1830 3633 -1710
rect -18500 -2297 3633 -1830
rect 4287 -1710 15673 -1703
rect 4287 -1830 5857 -1710
rect 5977 -1830 6857 -1710
rect 6977 -1830 15673 -1710
rect 4287 -2297 15673 -1830
rect 16327 -1710 38390 -1703
rect 16327 -1830 20260 -1710
rect 20380 -1830 22260 -1710
rect 22380 -1830 24260 -1710
rect 24380 -1830 26260 -1710
rect 26380 -1830 28260 -1710
rect 28380 -1830 30260 -1710
rect 30380 -1830 32260 -1710
rect 32380 -1830 34260 -1710
rect 34380 -1830 36260 -1710
rect 36380 -1830 38260 -1710
rect 38380 -1830 38390 -1710
rect 16327 -2297 38390 -1830
rect -18500 -2300 38390 -2297
rect 9000 -2600 11000 -2300
<< via4 >>
rect 40100 712 40220 832
rect -18900 -380 -18300 -80
rect -16900 -380 -16300 -80
rect -14900 -380 -14300 -80
rect -12900 -380 -12300 -80
rect -10900 -380 -10300 -80
rect -8900 -380 -8300 -80
rect -6900 -380 -6300 -80
rect -4900 -380 -4300 -80
rect -2900 -380 -2300 -80
rect -900 -380 -300 -80
rect 20260 -380 20860 -80
rect 22260 -380 22860 -80
rect 24260 -380 24860 -80
rect 26260 -380 26860 -80
rect 28260 -380 28860 -80
rect 30260 -380 30860 -80
rect 32260 -380 32860 -80
rect 34260 -380 34860 -80
rect 36260 -380 36860 -80
rect 38260 -380 38860 -80
rect -20480 -1480 -20120 -520
rect 40080 -1480 40440 -520
<< metal5 >>
rect -20500 45200 -300 45600
rect -20500 -520 -20100 45200
rect -18900 45000 -18300 45200
rect -16900 45000 -16300 45200
rect -14900 45000 -14300 45200
rect -12900 45000 -12300 45200
rect -10900 45000 -10300 45200
rect -8900 45000 -8300 45200
rect -6900 45000 -6300 45200
rect -4900 45000 -4300 45200
rect -2900 45000 -2300 45200
rect -900 45000 -300 45200
rect 20260 45200 40460 45600
rect 20260 45000 20860 45200
rect 22260 45000 22860 45200
rect 24260 45000 24860 45200
rect 26260 45000 26860 45200
rect 28260 45000 28860 45200
rect 30260 45000 30860 45200
rect 32260 45000 32860 45200
rect 34260 45000 34860 45200
rect 36260 45000 36860 45200
rect 38260 45000 38860 45200
rect 40060 832 40460 45200
rect 40060 712 40100 832
rect 40220 712 40460 832
rect -20500 -1480 -20480 -520
rect -20120 -1480 -20100 -520
rect -19900 -600 -19300 0
rect -18900 -60 -18300 0
rect -18920 -80 -18280 -60
rect -18920 -380 -18900 -80
rect -18300 -380 -18280 -80
rect -18920 -400 -18280 -380
rect -17900 -600 -17300 0
rect -16900 -60 -16300 0
rect -16920 -80 -16280 -60
rect -16920 -380 -16900 -80
rect -16300 -380 -16280 -80
rect -16920 -400 -16280 -380
rect -15900 -600 -15300 0
rect -14900 -60 -14300 0
rect -14920 -80 -14280 -60
rect -14920 -380 -14900 -80
rect -14300 -380 -14280 -80
rect -14920 -400 -14280 -380
rect -13900 -600 -13300 0
rect -12900 -60 -12300 0
rect -12920 -80 -12280 -60
rect -12920 -380 -12900 -80
rect -12300 -380 -12280 -80
rect -12920 -400 -12280 -380
rect -11900 -600 -11300 0
rect -10900 -60 -10300 0
rect -10920 -80 -10280 -60
rect -10920 -380 -10900 -80
rect -10300 -380 -10280 -80
rect -10920 -400 -10280 -380
rect -9900 -600 -9300 0
rect -8900 -60 -8300 0
rect -8920 -80 -8280 -60
rect -8920 -380 -8900 -80
rect -8300 -380 -8280 -80
rect -8920 -400 -8280 -380
rect -7900 -600 -7300 0
rect -6900 -60 -6300 0
rect -6920 -80 -6280 -60
rect -6920 -380 -6900 -80
rect -6300 -380 -6280 -80
rect -6920 -400 -6280 -380
rect -5900 -600 -5300 0
rect -4900 -60 -4300 0
rect -4920 -80 -4280 -60
rect -4920 -380 -4900 -80
rect -4300 -380 -4280 -80
rect -4920 -400 -4280 -380
rect -3900 -600 -3300 0
rect -2900 -60 -2300 0
rect -2920 -80 -2280 -60
rect -2920 -380 -2900 -80
rect -2300 -380 -2280 -80
rect -2920 -400 -2280 -380
rect -1900 -600 -1300 0
rect -900 -60 -300 0
rect 20260 -60 20860 0
rect -920 -80 -280 -60
rect -920 -380 -900 -80
rect -300 -380 -280 -80
rect -920 -400 -280 -380
rect 20240 -80 20880 -60
rect 20240 -380 20260 -80
rect 20860 -380 20880 -80
rect 20240 -400 20880 -380
rect 21260 -600 21860 0
rect 22260 -60 22860 0
rect 22240 -80 22880 -60
rect 22240 -380 22260 -80
rect 22860 -380 22880 -80
rect 22240 -400 22880 -380
rect 23260 -600 23860 0
rect 24260 -60 24860 0
rect 24240 -80 24880 -60
rect 24240 -380 24260 -80
rect 24860 -380 24880 -80
rect 24240 -400 24880 -380
rect 25260 -600 25860 0
rect 26260 -60 26860 0
rect 26240 -80 26880 -60
rect 26240 -380 26260 -80
rect 26860 -380 26880 -80
rect 26240 -400 26880 -380
rect 27260 -600 27860 0
rect 28260 -60 28860 0
rect 28240 -80 28880 -60
rect 28240 -380 28260 -80
rect 28860 -380 28880 -80
rect 28240 -400 28880 -380
rect 29260 -600 29860 0
rect 30260 -60 30860 0
rect 30240 -80 30880 -60
rect 30240 -380 30260 -80
rect 30860 -380 30880 -80
rect 30240 -400 30880 -380
rect 31260 -600 31860 0
rect 32260 -60 32860 0
rect 32240 -80 32880 -60
rect 32240 -380 32260 -80
rect 32860 -380 32880 -80
rect 32240 -400 32880 -380
rect 33260 -600 33860 0
rect 34260 -60 34860 0
rect 34240 -80 34880 -60
rect 34240 -380 34260 -80
rect 34860 -380 34880 -80
rect 34240 -400 34880 -380
rect 35260 -600 35860 0
rect 36260 -60 36860 0
rect 36240 -80 36880 -60
rect 36240 -380 36260 -80
rect 36860 -380 36880 -80
rect 36240 -400 36880 -380
rect 37260 -600 37860 0
rect 38260 -60 38860 0
rect 38240 -80 38880 -60
rect 38240 -380 38260 -80
rect 38860 -380 38880 -80
rect 38240 -400 38880 -380
rect 39260 -600 39860 0
rect -19900 -1400 39860 -600
rect 40060 -520 40460 712
rect -20500 -1500 -20100 -1480
rect 34400 -2600 36600 -1400
rect 40060 -1480 40080 -520
rect 40440 -1480 40460 -520
rect 40060 -1500 40460 -1480
use array_column_decode  array_column_decode_0
timestamp 1717569530
transform 0 1 -520 -1 0 3560
box -2020 6520 1560 13936
use array_core_block0  array_core_block0_0
timestamp 1717597427
transform 1 0 -20000 0 1 30696
box -33 -696 19983 14118
use array_core_block1  array_core_block1_0
timestamp 1717597427
transform 1 0 -20000 0 1 15000
box -33 0 19983 14814
use array_core_block2  array_core_block2_0
timestamp 1717597427
transform 1 0 -20000 0 1 0
box -33 0 19983 14819
use array_core_block3_alt  array_core_block3_alt_0
timestamp 1717597306
transform -1 0 39983 0 1 30000
box 0 0 19983 14623
use array_core_block4_alt  array_core_block4_alt_0
timestamp 1717597427
transform -1 0 39983 0 1 15000
box -33 0 19983 14623
use array_core_block5  array_core_block5_0
timestamp 1717597427
transform -1 0 39983 0 1 0
box -33 0 19983 14623
use array_core_block_routing  array_core_block_routing_0
array 0 0 -20040 0 2 15000
timestamp 1717570868
transform -1 0 40760 0 1 0
box 800 0 20840 15000
use array_core_block_routing  array_core_block_routing_1
array 0 0 19760 0 2 15000
timestamp 1717570868
transform 1 0 -20800 0 1 0
box 800 0 20840 15000
use array_row_decode  array_row_decode_0
timestamp 1717570567
transform 1 0 13210 0 1 28832
box -2020 168 1560 14074
use array_row_decode  array_row_decode_1
timestamp 1717570567
transform -1 0 6750 0 1 28832
box -2020 168 1560 14074
use lsi1v8o5v0  lsi1v8o5v0_0
array 0 0 1161 0 31 -400
timestamp 1717570567
transform -1 0 5048 0 -1 29307
box -42 -60 1371 293
use lsi1v8o5v0  lsi1v8o5v0_1
array 0 0 1161 0 31 -400
timestamp 1717570567
transform 1 0 14912 0 -1 29307
box -42 -60 1371 293
use lsi1v8o5v0  lsi1v8o5v0_2
array 0 0 1161 0 15 -400
timestamp 1717570567
transform 0 -1 6355 -1 0 1858
box -42 -60 1371 293
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1717569530
transform 1 0 15400 0 1 19900
box 0 0 1141 1169
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield_1
timestamp 1717569530
transform 1 0 3300 0 1 19900
box 0 0 1141 1169
use tg5v0  tg5v0_0
array 0 0 -800 0 9 2000
timestamp 1717597221
transform 0 -1 90 -1 0 -983
box 14 0 817 445
use tg5v0  tg5v0_1
array 0 0 -800 0 9 2000
timestamp 1717597221
transform 0 1 19869 -1 0 -983
box 14 0 817 445
use tg5v0  tg5v0_2
timestamp 1717597221
transform 0 -1 7385 -1 0 -983
box 14 0 817 445
use tg5v0  tg5v0_3
timestamp 1717597221
transform 0 -1 1385 -1 0 -983
box 14 0 817 445
use tg5v0  tg5v0_4
timestamp 1717597221
transform 0 -1 6385 -1 0 -983
box 14 0 817 445
use vb_divider  vb_divider_0
timestamp 1717569530
transform -1 0 11259 0 1 18400
box 0 0 759 986
<< labels >>
flabel metal2 8770 42772 11190 42872 0 FreeSans 320 0 0 0 a[8]
flabel metal2 8770 42634 11190 42734 0 FreeSans 320 0 0 0 a[7]
flabel metal2 8770 42496 11190 42596 0 FreeSans 320 0 0 0 a[6]
flabel metal2 8770 42358 11190 42458 0 FreeSans 320 0 0 0 a[5]
flabel metal2 8770 42220 11190 42320 0 FreeSans 320 0 0 0 a[4]
flabel metal3 8774 42880 8974 42960 0 FreeSans 320 0 0 0 a[0]
flabel metal3 9042 42880 9242 42960 0 FreeSans 320 0 0 0 a[1]
flabel metal3 9310 42880 9510 42960 0 FreeSans 320 0 0 0 a[2]
flabel metal3 9578 42880 9778 42960 0 FreeSans 320 0 0 0 a[3]
flabel metal3 10114 42880 10314 42960 0 FreeSans 320 0 0 0 a[5]
flabel metal3 10382 42880 10582 42960 0 FreeSans 320 0 0 0 a[6]
flabel metal3 10650 42880 10850 42960 0 FreeSans 320 0 0 0 a[7]
flabel metal3 10918 42880 11118 42960 0 FreeSans 320 0 0 0 a[8]
flabel metal3 9846 42880 10046 42960 0 FreeSans 320 0 0 0 a[4]
flabel metal2 4989 41532 5047 41590 0 FreeSans 160 0 0 0 l_w[0]
flabel metal2 4989 41132 5047 41190 0 FreeSans 160 0 0 0 l_w[1]
flabel metal2 4989 40732 5047 40790 0 FreeSans 160 0 0 0 l_w[2]
flabel metal2 4989 40332 5047 40390 0 FreeSans 160 0 0 0 l_w[3]
flabel metal2 4989 39932 5047 39990 0 FreeSans 160 0 0 0 l_w[4]
flabel metal2 4989 39532 5047 39590 0 FreeSans 160 0 0 0 l_w[5]
flabel metal2 4989 39132 5047 39190 0 FreeSans 160 0 0 0 l_w[6]
flabel metal2 4989 38732 5047 38790 0 FreeSans 160 0 0 0 l_w[7]
flabel metal2 4989 38332 5047 38390 0 FreeSans 160 0 0 0 l_w[8]
flabel metal2 4989 37932 5047 37990 0 FreeSans 160 0 0 0 l_w[9]
flabel metal2 4989 37532 5047 37590 0 FreeSans 160 0 0 0 l_w[10]
flabel metal2 4989 37132 5047 37190 0 FreeSans 160 0 0 0 l_w[11]
flabel metal2 4989 36732 5047 36790 0 FreeSans 160 0 0 0 l_w[12]
flabel metal2 4989 36332 5047 36390 0 FreeSans 160 0 0 0 l_w[13]
flabel metal2 4989 35932 5047 35990 0 FreeSans 160 0 0 0 l_w[14]
flabel metal2 4989 35532 5047 35590 0 FreeSans 160 0 0 0 l_w[15]
flabel metal2 4989 35132 5047 35190 0 FreeSans 160 0 0 0 l_w[16]
flabel metal2 4989 34732 5047 34790 0 FreeSans 160 0 0 0 l_w[17]
flabel metal2 4989 34332 5047 34390 0 FreeSans 160 0 0 0 l_w[18]
flabel metal2 4989 33932 5047 33990 0 FreeSans 160 0 0 0 l_w[19]
flabel metal2 4989 33532 5047 33590 0 FreeSans 160 0 0 0 l_w[20]
flabel metal2 4989 33132 5047 33190 0 FreeSans 160 0 0 0 l_w[21]
flabel metal2 4989 32732 5047 32790 0 FreeSans 160 0 0 0 l_w[22]
flabel metal2 4989 32332 5047 32390 0 FreeSans 160 0 0 0 l_w[23]
flabel metal2 4989 31932 5047 31990 0 FreeSans 160 0 0 0 l_w[24]
flabel metal2 4989 31532 5047 31590 0 FreeSans 160 0 0 0 l_w[25]
flabel metal2 4989 31132 5047 31190 0 FreeSans 160 0 0 0 l_w[26]
flabel metal2 4989 30732 5047 30790 0 FreeSans 160 0 0 0 l_w[27]
flabel metal2 4989 30332 5047 30390 0 FreeSans 160 0 0 0 l_w[28]
flabel metal2 4989 29932 5047 29990 0 FreeSans 160 0 0 0 l_w[29]
flabel metal2 4989 29532 5047 29590 0 FreeSans 160 0 0 0 l_w[30]
flabel metal2 4989 29132 5047 29190 0 FreeSans 160 0 0 0 l_w[31]
flabel metal2 14913 41532 14971 41590 0 FreeSans 160 0 0 0 r_w[0]
flabel metal2 14913 41132 14971 41190 0 FreeSans 160 0 0 0 r_w[1]
flabel metal2 14913 40732 14971 40790 0 FreeSans 160 0 0 0 r_w[2]
flabel metal2 14913 40332 14971 40390 0 FreeSans 160 0 0 0 r_w[3]
flabel metal2 14913 39932 14971 39990 0 FreeSans 160 0 0 0 r_w[4]
flabel metal2 14913 39532 14971 39590 0 FreeSans 160 0 0 0 r_w[5]
flabel metal2 14913 39132 14971 39190 0 FreeSans 160 0 0 0 r_w[6]
flabel metal2 14913 38732 14971 38790 0 FreeSans 160 0 0 0 r_w[7]
flabel metal2 14913 38332 14971 38390 0 FreeSans 160 0 0 0 r_w[8]
flabel metal2 14913 37932 14971 37990 0 FreeSans 160 0 0 0 r_w[9]
flabel metal2 14913 37532 14971 37590 0 FreeSans 160 0 0 0 r_w[10]
flabel metal2 14913 37132 14971 37190 0 FreeSans 160 0 0 0 r_w[11]
flabel metal2 14913 36732 14971 36790 0 FreeSans 160 0 0 0 r_w[12]
flabel metal2 14913 36332 14971 36390 0 FreeSans 160 0 0 0 r_w[13]
flabel metal2 14913 35932 14971 35990 0 FreeSans 160 0 0 0 r_w[14]
flabel metal2 14913 35532 14971 35590 0 FreeSans 160 0 0 0 r_w[15]
flabel metal2 14913 35132 14971 35190 0 FreeSans 160 0 0 0 r_w[16]
flabel metal2 14913 34732 14971 34790 0 FreeSans 160 0 0 0 r_w[17]
flabel metal2 14913 34332 14971 34390 0 FreeSans 160 0 0 0 r_w[18]
flabel metal2 14913 33932 14971 33990 0 FreeSans 160 0 0 0 r_w[19]
flabel metal2 14913 33532 14971 33590 0 FreeSans 160 0 0 0 r_w[20]
flabel metal2 14913 33132 14971 33190 0 FreeSans 160 0 0 0 r_w[21]
flabel metal2 14913 32732 14971 32790 0 FreeSans 160 0 0 0 r_w[22]
flabel metal2 14913 32332 14971 32390 0 FreeSans 160 0 0 0 r_w[23]
flabel metal2 14913 31932 14971 31990 0 FreeSans 160 0 0 0 r_w[24]
flabel metal2 14913 31532 14971 31590 0 FreeSans 160 0 0 0 r_w[25]
flabel metal2 14913 31132 14971 31190 0 FreeSans 160 0 0 0 r_w[26]
flabel metal2 14913 30732 14971 30790 0 FreeSans 160 0 0 0 r_w[27]
flabel metal2 14913 30332 14971 30390 0 FreeSans 160 0 0 0 r_w[28]
flabel metal2 14913 29932 14971 29990 0 FreeSans 160 0 0 0 r_w[29]
flabel metal2 14913 29532 14971 29590 0 FreeSans 160 0 0 0 r_w[30]
flabel metal2 14913 29132 14971 29190 0 FreeSans 160 0 0 0 r_w[31]
flabel metal5 -19900 -1400 38500 -600 0 FreeSans 3200 0 0 0 VTUN
flabel metal4 40 400 540 44300 0 FreeSans 800 0 0 0 VINJ
flabel metal3 40 230 440 43820 0 FreeSans 1600 0 0 0 vb
flabel metal2 12180 1799 12238 1857 0 FreeSans 160 0 0 0 c[0]
flabel metal2 11780 1799 11838 1857 0 FreeSans 160 0 0 0 c[1]
flabel metal2 11380 1799 11438 1857 0 FreeSans 160 0 0 0 c[2]
flabel metal2 10980 1799 11038 1857 0 FreeSans 160 0 0 0 c[3]
flabel metal2 10580 1799 10638 1857 0 FreeSans 160 0 0 0 c[4]
flabel metal2 10180 1799 10238 1857 0 FreeSans 160 0 0 0 c[5]
flabel metal2 9780 1799 9838 1857 0 FreeSans 160 0 0 0 c[6]
flabel metal2 9380 1799 9438 1857 0 FreeSans 160 0 0 0 c[7]
flabel metal2 8980 1799 9038 1857 0 FreeSans 160 0 0 0 c[8]
flabel metal2 8580 1799 8638 1857 0 FreeSans 160 0 0 0 c[9]
flabel metal2 8180 1799 8238 1857 0 FreeSans 160 0 0 0 c[10]
flabel metal2 7780 1799 7838 1857 0 FreeSans 160 0 0 0 c[11]
flabel metal2 7380 1799 7438 1857 0 FreeSans 160 0 0 0 c[12]
flabel metal2 6980 1799 7038 1857 0 FreeSans 160 0 0 0 c[13]
flabel metal2 6580 1799 6638 1857 0 FreeSans 160 0 0 0 c[14]
flabel metal2 6180 1799 6238 1857 0 FreeSans 160 0 0 0 c[15]
flabel metal3 4600 4400 4800 4600 0 FreeSans 800 0 0 0 VPWR
flabel metal3 15100 4400 15300 4600 0 FreeSans 800 0 0 0 VPWR
flabel metal3 14300 4400 14500 4600 0 FreeSans 800 0 0 0 VGND
flabel metal3 5400 4400 5600 4600 0 FreeSans 800 0 0 0 VGND
flabel metal3 3800 4400 4000 4600 0 FreeSans 800 0 0 0 vinj
flabel metal3 15900 4400 16100 4600 0 FreeSans 800 0 0 0 vinj
flabel metal4 3630 -2300 16330 -1700 0 FreeSans 3200 0 0 0 VINJ
flabel metal1 -110 -2200 90 -2000 0 FreeSans 400 0 0 0 l_vout
flabel metal3 -18600 -600 800 -200 0 FreeSans 800 0 0 0 VSRC
flabel metal3 3000 4400 3200 4600 0 FreeSans 800 0 0 0 VCTRL
flabel pwell 3333 19933 4408 21036 0 FreeSans 160 0 0 0 VGND
flabel metal1 3300 21069 4441 21090 0 FreeSans 160 0 0 0 VGND
flabel pwell 15433 19933 16508 21036 0 FreeSans 160 0 0 0 VGND
flabel metal1 15444 21069 16541 21090 0 FreeSans 160 0 0 0 VGND
flabel metal4 -18900 -1500 33776 -500 0 FreeSans 3200 0 0 0 VGND
flabel metal3 7300 45500 7500 45600 0 FreeSans 400 0 0 0 a[0]
port 3 nsew
flabel metal3 7900 45500 8100 45600 0 FreeSans 400 0 0 0 a[1]
port 4 nsew signal input
flabel metal3 8500 45500 8700 45600 0 FreeSans 400 0 0 0 a[2]
port 5 nsew signal input
flabel metal3 9100 45500 9300 45600 0 FreeSans 400 0 0 0 a[3]
port 6 nsew signal input
flabel metal3 9700 45500 9900 45600 0 FreeSans 400 0 0 0 a[4]
port 7 nsew signal input
flabel metal3 10300 45500 10500 45600 0 FreeSans 400 0 0 0 a[5]
port 8 nsew signal input
flabel metal3 10900 45500 11100 45600 0 FreeSans 400 0 0 0 a[6]
port 9 nsew signal input
flabel metal3 11500 45500 11700 45600 0 FreeSans 400 0 0 0 a[7]
port 10 nsew signal input
flabel metal3 12100 45500 12300 45600 0 FreeSans 400 0 0 0 a[8]
port 11 nsew signal input
flabel metal3 12700 45500 13500 45600 0 FreeSans 400 0 0 0 VPWR
port 1 nsew power default
flabel metal3 6100 45500 6900 45600 0 FreeSans 400 0 0 0 VGND
port 2 nsew ground default
flabel metal3 2860 -2600 3520 -2400 0 FreeSans 800 0 0 0 VCTRL
port 15 nsew
flabel metal3 2090 -2600 2750 -2400 0 FreeSans 800 0 0 0 VSRC
port 16 nsew
flabel metal4 9000 -2600 11000 -2400 0 FreeSans 800 0 0 0 VINJ
port 13 nsew
flabel metal3 4400 -2600 4800 -2400 0 FreeSans 800 0 0 0 VOUT0
port 14 nsew
flabel metal5 34400 -2600 36600 -2400 0 FreeSans 1600 0 0 0 VTUN
port 12 nsew
flabel metal3 23900 -2600 26100 -2400 0 FreeSans 1600 0 0 0 VGND
port 2 nsew
flabel metal4 100 -400 19400 100 0 FreeSans 1600 0 0 0 VSRC
flabel metal2 3677 29131 3727 29181 0 FreeSans 80 0 0 0 l_row_en_b[31]
flabel metal2 3677 29531 3727 29581 0 FreeSans 80 0 0 0 l_row_en_b[30]
flabel metal2 3677 29931 3727 29981 0 FreeSans 80 0 0 0 l_row_en_b[29]
flabel metal2 3677 30331 3727 30381 0 FreeSans 80 0 0 0 l_row_en_b[28]
flabel metal2 3677 30731 3727 30781 0 FreeSans 80 0 0 0 l_row_en_b[27]
flabel metal2 3677 31131 3727 31181 0 FreeSans 80 0 0 0 l_row_en_b[26]
flabel metal2 3677 31531 3727 31581 0 FreeSans 80 0 0 0 l_row_en_b[25]
flabel metal2 3677 31931 3727 31981 0 FreeSans 80 0 0 0 l_row_en_b[24]
flabel metal2 3677 32331 3727 32381 0 FreeSans 80 0 0 0 l_row_en_b[23]
flabel metal2 3677 32731 3727 32781 0 FreeSans 80 0 0 0 l_row_en_b[22]
flabel metal2 3677 33131 3727 33181 0 FreeSans 80 0 0 0 l_row_en_b[21]
flabel metal2 3677 33531 3727 33581 0 FreeSans 80 0 0 0 l_row_en_b[20]
flabel metal2 3677 33931 3727 33981 0 FreeSans 80 0 0 0 l_row_en_b[19]
flabel metal2 3677 34331 3727 34381 0 FreeSans 80 0 0 0 l_row_en_b[18]
flabel metal2 3677 34731 3727 34781 0 FreeSans 80 0 0 0 l_row_en_b[17]
flabel metal2 3677 35131 3727 35181 0 FreeSans 80 0 0 0 l_row_en_b[16]
flabel metal2 3677 35531 3727 35581 0 FreeSans 80 0 0 0 l_row_en_b[15]
flabel metal2 3677 35931 3727 35981 0 FreeSans 80 0 0 0 l_row_en_b[14]
flabel metal2 3677 36331 3727 36381 0 FreeSans 80 0 0 0 l_row_en_b[13]
flabel metal2 3677 36731 3727 36781 0 FreeSans 80 0 0 0 l_row_en_b[12]
flabel metal2 3677 37131 3727 37181 0 FreeSans 80 0 0 0 l_row_en_b[11]
flabel metal2 3677 37531 3727 37581 0 FreeSans 80 0 0 0 l_row_en_b[10]
flabel metal2 3677 37931 3727 37981 0 FreeSans 80 0 0 0 l_row_en_b[9]
flabel metal2 3677 38331 3727 38381 0 FreeSans 80 0 0 0 l_row_en_b[8]
flabel metal2 3677 38731 3727 38781 0 FreeSans 80 0 0 0 l_row_en_b[7]
flabel metal2 3677 39131 3727 39181 0 FreeSans 80 0 0 0 l_row_en_b[6]
flabel metal2 3677 39531 3727 39581 0 FreeSans 80 0 0 0 l_row_en_b[5]
flabel metal2 3677 39931 3727 39981 0 FreeSans 80 0 0 0 l_row_en_b[4]
flabel metal2 3677 40331 3727 40381 0 FreeSans 80 0 0 0 l_row_en_b[3]
flabel metal2 3677 40731 3727 40781 0 FreeSans 80 0 0 0 l_row_en_b[2]
flabel metal2 3677 41131 3727 41181 0 FreeSans 80 0 0 0 l_row_en_b[1]
flabel metal2 3677 41531 3727 41581 0 FreeSans 80 0 0 0 l_row_en_b[0]
flabel metal2 3677 29195 3727 29245 0 FreeSans 80 0 0 0 l_row_en[31]
flabel metal2 3677 29595 3727 29645 0 FreeSans 80 0 0 0 l_row_en[30]
flabel metal2 3677 29995 3727 30045 0 FreeSans 80 0 0 0 l_row_en[29]
flabel metal2 3677 30395 3727 30445 0 FreeSans 80 0 0 0 l_row_en[28]
flabel metal2 3677 30795 3727 30845 0 FreeSans 80 0 0 0 l_row_en[27]
flabel metal2 3677 31195 3727 31245 0 FreeSans 80 0 0 0 l_row_en[26]
flabel metal2 3677 31595 3727 31645 0 FreeSans 80 0 0 0 l_row_en[25]
flabel metal2 3677 31995 3727 32045 0 FreeSans 80 0 0 0 l_row_en[24]
flabel metal2 3677 32395 3727 32445 0 FreeSans 80 0 0 0 l_row_en[23]
flabel metal2 3677 32795 3727 32845 0 FreeSans 80 0 0 0 l_row_en[22]
flabel metal2 3677 33195 3727 33245 0 FreeSans 80 0 0 0 l_row_en[21]
flabel metal2 3677 33595 3727 33645 0 FreeSans 80 0 0 0 l_row_en[20]
flabel metal2 3677 33995 3727 34045 0 FreeSans 80 0 0 0 l_row_en[19]
flabel metal2 3677 34395 3727 34445 0 FreeSans 80 0 0 0 l_row_en[18]
flabel metal2 3677 34795 3727 34845 0 FreeSans 80 0 0 0 l_row_en[17]
flabel metal2 3677 35195 3727 35245 0 FreeSans 80 0 0 0 l_row_en[16]
flabel metal2 3677 35595 3727 35645 0 FreeSans 80 0 0 0 l_row_en[15]
flabel metal2 3677 35995 3727 36045 0 FreeSans 80 0 0 0 l_row_en[14]
flabel metal2 3677 36395 3727 36445 0 FreeSans 80 0 0 0 l_row_en[13]
flabel metal2 3677 36795 3727 36845 0 FreeSans 80 0 0 0 l_row_en[12]
flabel metal2 3677 37195 3727 37245 0 FreeSans 80 0 0 0 l_row_en[11]
flabel metal2 3677 37595 3727 37645 0 FreeSans 80 0 0 0 l_row_en[10]
flabel metal2 3677 37995 3727 38045 0 FreeSans 80 0 0 0 l_row_en[9]
flabel metal2 3677 38395 3727 38445 0 FreeSans 80 0 0 0 l_row_en[8]
flabel metal2 3677 38795 3727 38845 0 FreeSans 80 0 0 0 l_row_en[7]
flabel metal2 3677 39195 3727 39245 0 FreeSans 80 0 0 0 l_row_en[6]
flabel metal2 3677 39595 3727 39645 0 FreeSans 80 0 0 0 l_row_en[5]
flabel metal2 3677 39995 3727 40045 0 FreeSans 80 0 0 0 l_row_en[4]
flabel metal2 3677 40395 3727 40445 0 FreeSans 80 0 0 0 l_row_en[3]
flabel metal2 3677 40795 3727 40845 0 FreeSans 80 0 0 0 l_row_en[2]
flabel metal2 3677 41195 3727 41245 0 FreeSans 80 0 0 0 l_row_en[1]
flabel metal2 3677 41595 3727 41645 0 FreeSans 80 0 0 0 l_row_en[0]
flabel metal2 16233 29131 16283 29181 0 FreeSans 80 0 0 0 r_row_en_b[31]
flabel metal2 16233 29531 16283 29581 0 FreeSans 80 0 0 0 r_row_en_b[30]
flabel metal2 16233 29931 16283 29981 0 FreeSans 80 0 0 0 r_row_en_b[29]
flabel metal2 16233 30331 16283 30381 0 FreeSans 80 0 0 0 r_row_en_b[28]
flabel metal2 16233 30731 16283 30781 0 FreeSans 80 0 0 0 r_row_en_b[27]
flabel metal2 16233 31131 16283 31181 0 FreeSans 80 0 0 0 r_row_en_b[26]
flabel metal2 16233 31531 16283 31581 0 FreeSans 80 0 0 0 r_row_en_b[25]
flabel metal2 16233 31931 16283 31981 0 FreeSans 80 0 0 0 r_row_en_b[24]
flabel metal2 16233 32331 16283 32381 0 FreeSans 80 0 0 0 r_row_en_b[23]
flabel metal2 16233 32731 16283 32781 0 FreeSans 80 0 0 0 r_row_en_b[22]
flabel metal2 16233 33131 16283 33181 0 FreeSans 80 0 0 0 r_row_en_b[21]
flabel metal2 16233 33531 16283 33581 0 FreeSans 80 0 0 0 r_row_en_b[20]
flabel metal2 16233 33931 16283 33981 0 FreeSans 80 0 0 0 r_row_en_b[19]
flabel metal2 16233 34331 16283 34381 0 FreeSans 80 0 0 0 r_row_en_b[18]
flabel metal2 16233 34731 16283 34781 0 FreeSans 80 0 0 0 r_row_en_b[17]
flabel metal2 16233 35131 16283 35181 0 FreeSans 80 0 0 0 r_row_en_b[16]
flabel metal2 16233 35531 16283 35581 0 FreeSans 80 0 0 0 r_row_en_b[15]
flabel metal2 16233 35931 16283 35981 0 FreeSans 80 0 0 0 r_row_en_b[14]
flabel metal2 16233 36331 16283 36381 0 FreeSans 80 0 0 0 r_row_en_b[13]
flabel metal2 16233 36731 16283 36781 0 FreeSans 80 0 0 0 r_row_en_b[12]
flabel metal2 16233 37131 16283 37181 0 FreeSans 80 0 0 0 r_row_en_b[11]
flabel metal2 16233 37531 16283 37581 0 FreeSans 80 0 0 0 r_row_en_b[10]
flabel metal2 16233 37931 16283 37981 0 FreeSans 80 0 0 0 r_row_en_b[9]
flabel metal2 16233 38331 16283 38381 0 FreeSans 80 0 0 0 r_row_en_b[8]
flabel metal2 16233 38731 16283 38781 0 FreeSans 80 0 0 0 r_row_en_b[7]
flabel metal2 16233 39131 16283 39181 0 FreeSans 80 0 0 0 r_row_en_b[6]
flabel metal2 16233 39531 16283 39581 0 FreeSans 80 0 0 0 r_row_en_b[5]
flabel metal2 16233 39931 16283 39981 0 FreeSans 80 0 0 0 r_row_en_b[4]
flabel metal2 16233 40331 16283 40381 0 FreeSans 80 0 0 0 r_row_en_b[3]
flabel metal2 16233 40731 16283 40781 0 FreeSans 80 0 0 0 r_row_en_b[2]
flabel metal2 16233 41131 16283 41181 0 FreeSans 80 0 0 0 r_row_en_b[1]
flabel metal2 16233 41531 16283 41581 0 FreeSans 80 0 0 0 r_row_en_b[0]
flabel metal2 16233 29195 16283 29245 0 FreeSans 80 0 0 0 r_row_en[31]
flabel metal2 16233 29595 16283 29645 0 FreeSans 80 0 0 0 r_row_en[30]
flabel metal2 16233 29995 16283 30045 0 FreeSans 80 0 0 0 r_row_en[29]
flabel metal2 16233 30395 16283 30445 0 FreeSans 80 0 0 0 r_row_en[28]
flabel metal2 16233 30795 16283 30845 0 FreeSans 80 0 0 0 r_row_en[27]
flabel metal2 16233 31195 16283 31245 0 FreeSans 80 0 0 0 r_row_en[26]
flabel metal2 16233 31595 16283 31645 0 FreeSans 80 0 0 0 r_row_en[25]
flabel metal2 16233 31995 16283 32045 0 FreeSans 80 0 0 0 r_row_en[24]
flabel metal2 16233 32395 16283 32445 0 FreeSans 80 0 0 0 r_row_en[23]
flabel metal2 16233 32795 16283 32845 0 FreeSans 80 0 0 0 r_row_en[22]
flabel metal2 16233 33195 16283 33245 0 FreeSans 80 0 0 0 r_row_en[21]
flabel metal2 16233 33595 16283 33645 0 FreeSans 80 0 0 0 r_row_en[20]
flabel metal2 16233 33995 16283 34045 0 FreeSans 80 0 0 0 r_row_en[19]
flabel metal2 16233 34395 16283 34445 0 FreeSans 80 0 0 0 r_row_en[18]
flabel metal2 16233 34795 16283 34845 0 FreeSans 80 0 0 0 r_row_en[17]
flabel metal2 16233 35195 16283 35245 0 FreeSans 80 0 0 0 r_row_en[16]
flabel metal2 16233 35595 16283 35645 0 FreeSans 80 0 0 0 r_row_en[15]
flabel metal2 16233 35995 16283 36045 0 FreeSans 80 0 0 0 r_row_en[14]
flabel metal2 16233 36395 16283 36445 0 FreeSans 80 0 0 0 r_row_en[13]
flabel metal2 16233 36795 16283 36845 0 FreeSans 80 0 0 0 r_row_en[12]
flabel metal2 16233 37195 16283 37245 0 FreeSans 80 0 0 0 r_row_en[11]
flabel metal2 16233 37595 16283 37645 0 FreeSans 80 0 0 0 r_row_en[10]
flabel metal2 16233 37995 16283 38045 0 FreeSans 80 0 0 0 r_row_en[9]
flabel metal2 16233 38395 16283 38445 0 FreeSans 80 0 0 0 r_row_en[8]
flabel metal2 16233 38795 16283 38845 0 FreeSans 80 0 0 0 r_row_en[7]
flabel metal2 16233 39195 16283 39245 0 FreeSans 80 0 0 0 r_row_en[6]
flabel metal2 16233 39595 16283 39645 0 FreeSans 80 0 0 0 r_row_en[5]
flabel metal2 16233 39995 16283 40045 0 FreeSans 80 0 0 0 r_row_en[4]
flabel metal2 16233 40395 16283 40445 0 FreeSans 80 0 0 0 r_row_en[3]
flabel metal2 16233 40795 16283 40845 0 FreeSans 80 0 0 0 r_row_en[2]
flabel metal2 16233 41195 16283 41245 0 FreeSans 80 0 0 0 r_row_en[1]
flabel metal2 16233 41595 16283 41645 0 FreeSans 80 0 0 0 r_row_en[0]
flabel metal3 4100 45500 4900 45600 0 FreeSans 400 0 0 0 VPWR
port 1 nsew power default
flabel metal3 14700 45500 15500 45600 0 FreeSans 400 0 0 0 VGND
port 2 nsew ground default
flabel metal1 19400 -2200 19600 -2000 0 FreeSans 800 0 0 0 r_vout
flabel metal3 17200 -2600 17800 -2400 0 FreeSans 800 0 0 0 VOUT1
flabel metal3 19520 230 19920 43820 0 FreeSans 1600 0 0 0 vb
flabel metal4 19420 400 19920 44300 0 FreeSans 320 0 0 0 vinj
<< end >>
