magic
tech sky130A
magscale 1 2
timestamp 1717349067
<< polycont >>
rect 1524 -2400 1586 -2342
<< locali >>
rect 1502 -2331 1610 -2322
rect 1502 -2409 1516 -2331
rect 1594 -2409 1610 -2331
rect 1502 -2416 1610 -2409
<< viali >>
rect 1516 -2342 1594 -2331
rect 1516 -2400 1524 -2342
rect 1524 -2400 1586 -2342
rect 1586 -2400 1594 -2342
rect 1516 -2409 1594 -2400
<< metal1 >>
rect 1500 -2325 1610 -2320
rect 1500 -2415 1510 -2325
rect 1600 -2415 1610 -2325
rect 1500 -2420 1610 -2415
<< via1 >>
rect 1660 -2020 1730 -1960
rect 1510 -2331 1600 -2325
rect 1510 -2409 1516 -2331
rect 1516 -2409 1594 -2331
rect 1594 -2409 1600 -2331
rect 1510 -2415 1600 -2409
<< metal2 >>
rect 1650 -1960 1740 -1954
rect 1650 -2020 1659 -1960
rect 1730 -2020 1740 -1960
rect 1650 -2028 1740 -2020
rect 1500 -2325 1610 -2320
rect 1500 -2415 1510 -2325
rect 1600 -2415 1610 -2325
rect 1500 -2420 1610 -2415
<< via2 >>
rect 1659 -2020 1660 -1960
rect 1660 -2020 1730 -1960
rect 1515 -2410 1595 -2330
<< metal3 >>
rect 1470 -1830 1740 -1570
rect 1650 -1960 1740 -1830
rect 1650 -2020 1659 -1960
rect 1730 -2020 1740 -1960
rect 1650 -2030 1740 -2020
rect 1510 -2326 1600 -2320
rect 1505 -2414 1511 -2326
rect 1599 -2414 1605 -2326
rect 1510 -2420 1600 -2414
<< via3 >>
rect 1511 -2330 1599 -2326
rect 1511 -2410 1515 -2330
rect 1515 -2410 1595 -2330
rect 1595 -2410 1599 -2330
rect 1511 -2414 1599 -2410
<< mimcap >>
rect 1500 -1710 1700 -1600
rect 1500 -1780 1520 -1710
rect 1590 -1780 1700 -1710
rect 1500 -1800 1700 -1780
<< mimcapcontact >>
rect 1520 -1780 1590 -1710
<< metal4 >>
rect 1510 -1710 1600 -1700
rect 1510 -1780 1520 -1710
rect 1590 -1780 1600 -1710
rect 1510 -2326 1600 -1780
rect 1510 -2414 1511 -2326
rect 1599 -2414 1600 -2326
rect 1510 -2420 1600 -2414
use fgcell_amp  x1
timestamp 1717349067
transform 1 0 384 0 1 3012
box 140 -7210 4106 -4964
<< end >>
