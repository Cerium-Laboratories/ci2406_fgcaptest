magic
tech sky130A
timestamp 1717165718
<< nwell >>
rect -42 133 1119 293
<< pwell >>
rect -14 -60 1091 55
<< mvnmos >>
rect 20 0 70 50
rect 99 0 149 50
rect 237 0 287 50
rect 316 0 366 50
rect 454 0 504 50
rect 533 0 583 50
rect 612 0 662 50
rect 691 0 741 50
rect 770 0 820 50
rect 849 0 899 50
rect 928 0 978 50
rect 1007 0 1057 50
<< mvpmos >>
rect 20 166 70 216
rect 99 166 149 216
rect 237 166 287 216
rect 316 166 366 216
rect 454 166 504 216
rect 533 166 583 216
rect 612 166 662 216
rect 691 166 741 216
rect 770 166 820 216
rect 849 166 899 216
rect 928 166 978 216
rect 1007 166 1057 216
<< mvndiff >>
rect -9 46 20 50
rect -9 4 -3 46
rect 14 4 20 46
rect -9 0 20 4
rect 70 46 99 50
rect 70 4 76 46
rect 93 4 99 46
rect 70 0 99 4
rect 149 46 178 50
rect 149 4 155 46
rect 172 4 178 46
rect 149 0 178 4
rect 208 46 237 50
rect 208 4 214 46
rect 231 4 237 46
rect 208 0 237 4
rect 287 46 316 50
rect 287 4 293 46
rect 310 4 316 46
rect 287 0 316 4
rect 366 46 395 50
rect 366 4 372 46
rect 389 4 395 46
rect 366 0 395 4
rect 425 46 454 50
rect 425 4 431 46
rect 448 4 454 46
rect 425 0 454 4
rect 504 46 533 50
rect 504 4 510 46
rect 527 4 533 46
rect 504 0 533 4
rect 583 46 612 50
rect 583 4 589 46
rect 606 4 612 46
rect 583 0 612 4
rect 662 46 691 50
rect 662 4 668 46
rect 685 4 691 46
rect 662 0 691 4
rect 741 46 770 50
rect 741 4 747 46
rect 764 4 770 46
rect 741 0 770 4
rect 820 46 849 50
rect 820 4 826 46
rect 843 4 849 46
rect 820 0 849 4
rect 899 46 928 50
rect 899 4 905 46
rect 922 4 928 46
rect 899 0 928 4
rect 978 46 1007 50
rect 978 4 984 46
rect 1001 4 1007 46
rect 978 0 1007 4
rect 1057 46 1086 50
rect 1057 4 1063 46
rect 1080 4 1086 46
rect 1057 0 1086 4
<< mvpdiff >>
rect -9 212 20 216
rect -9 170 -3 212
rect 14 170 20 212
rect -9 166 20 170
rect 70 212 99 216
rect 70 170 76 212
rect 93 170 99 212
rect 70 166 99 170
rect 149 212 178 216
rect 149 170 155 212
rect 172 170 178 212
rect 149 166 178 170
rect 208 212 237 216
rect 208 170 214 212
rect 231 170 237 212
rect 208 166 237 170
rect 287 212 316 216
rect 287 170 293 212
rect 310 170 316 212
rect 287 166 316 170
rect 366 212 395 216
rect 366 170 372 212
rect 389 170 395 212
rect 366 166 395 170
rect 425 212 454 216
rect 425 170 431 212
rect 448 170 454 212
rect 425 166 454 170
rect 504 212 533 216
rect 504 170 510 212
rect 527 170 533 212
rect 504 166 533 170
rect 583 212 612 216
rect 583 170 589 212
rect 606 170 612 212
rect 583 166 612 170
rect 662 212 691 216
rect 662 170 668 212
rect 685 170 691 212
rect 662 166 691 170
rect 741 212 770 216
rect 741 170 747 212
rect 764 170 770 212
rect 741 166 770 170
rect 820 212 849 216
rect 820 170 826 212
rect 843 170 849 212
rect 820 166 849 170
rect 899 212 928 216
rect 899 170 905 212
rect 922 170 928 212
rect 899 166 928 170
rect 978 212 1007 216
rect 978 170 984 212
rect 1001 170 1007 212
rect 978 166 1007 170
rect 1057 212 1086 216
rect 1057 170 1063 212
rect 1080 170 1086 212
rect 1057 166 1086 170
<< mvndiffc >>
rect -3 4 14 46
rect 76 4 93 46
rect 155 4 172 46
rect 214 4 231 46
rect 293 4 310 46
rect 372 4 389 46
rect 431 4 448 46
rect 510 4 527 46
rect 589 4 606 46
rect 668 4 685 46
rect 747 4 764 46
rect 826 4 843 46
rect 905 4 922 46
rect 984 4 1001 46
rect 1063 4 1080 46
<< mvpdiffc >>
rect -3 170 14 212
rect 76 170 93 212
rect 155 170 172 212
rect 214 170 231 212
rect 293 170 310 212
rect 372 170 389 212
rect 431 170 448 212
rect 510 170 527 212
rect 589 170 606 212
rect 668 170 685 212
rect 747 170 764 212
rect 826 170 843 212
rect 905 170 922 212
rect 984 170 1001 212
rect 1063 170 1080 212
<< mvpsubdiff >>
rect -3 -60 9 -43
rect 1068 -60 1080 -43
<< mvnsubdiff >>
rect -3 243 9 260
rect 1068 243 1080 260
<< mvpsubdiffcont >>
rect 9 -60 1068 -43
<< mvnsubdiffcont >>
rect 9 243 1068 260
<< poly >>
rect 20 216 70 229
rect 99 216 149 229
rect 237 216 287 229
rect 316 216 366 229
rect 454 216 504 229
rect 533 216 583 229
rect 612 216 662 229
rect 691 216 741 229
rect 770 216 820 229
rect 849 216 899 229
rect 928 216 978 229
rect 1007 216 1057 229
rect 20 140 70 166
rect 20 123 31 140
rect 59 123 70 140
rect 20 50 70 123
rect 99 97 149 166
rect 237 142 287 166
rect 237 125 248 142
rect 276 125 287 142
rect 237 120 287 125
rect 316 142 366 166
rect 316 125 327 142
rect 355 125 366 142
rect 316 120 366 125
rect 454 158 504 166
rect 533 158 583 166
rect 612 158 662 166
rect 691 158 741 166
rect 454 131 741 158
rect 99 80 110 97
rect 138 80 149 97
rect 454 114 465 131
rect 493 114 741 131
rect 454 112 741 114
rect 770 158 820 166
rect 849 158 899 166
rect 928 158 978 166
rect 1007 158 1057 166
rect 770 141 1057 158
rect 99 50 149 80
rect 237 91 287 96
rect 237 74 248 91
rect 276 74 287 91
rect 237 50 287 74
rect 316 91 366 96
rect 316 74 327 91
rect 355 74 366 91
rect 316 50 366 74
rect 454 58 583 112
rect 454 50 504 58
rect 533 50 583 58
rect 612 86 741 91
rect 612 69 628 86
rect 645 69 741 86
rect 612 58 741 69
rect 612 50 662 58
rect 691 50 741 58
rect 770 75 775 141
rect 809 112 1057 141
rect 809 75 899 112
rect 770 58 899 75
rect 770 50 820 58
rect 849 50 899 58
rect 928 86 1057 91
rect 928 69 944 86
rect 961 69 1057 86
rect 928 58 1057 69
rect 928 50 978 58
rect 1007 50 1057 58
rect 20 -13 70 0
rect 99 -13 149 0
rect 237 -13 287 0
rect 316 -13 366 0
rect 454 -13 504 0
rect 533 -13 583 0
rect 612 -13 662 0
rect 691 -13 741 0
rect 770 -13 820 0
rect 849 -13 899 0
rect 928 -13 978 0
rect 1007 -13 1057 0
<< polycont >>
rect 31 123 59 140
rect 248 125 276 142
rect 327 125 355 142
rect 110 80 138 97
rect 465 114 493 131
rect 248 74 276 91
rect 327 74 355 91
rect 628 69 645 86
rect 775 75 809 141
rect 944 69 961 86
<< locali >>
rect -3 243 9 260
rect 1068 254 1080 260
rect -3 212 14 220
rect -3 97 14 170
rect 76 212 93 220
rect 76 162 93 170
rect 155 212 172 220
rect 31 140 59 148
rect 31 115 59 123
rect -3 46 14 80
rect 110 97 138 105
rect 110 72 138 80
rect 155 57 172 170
rect -3 -4 14 4
rect 76 46 93 54
rect 76 -21 93 4
rect 155 -4 172 4
rect 214 212 231 220
rect 293 212 310 237
rect 293 162 310 170
rect 372 212 389 220
rect 214 46 231 159
rect 248 142 276 150
rect 248 117 276 125
rect 327 148 332 165
rect 350 148 355 165
rect 327 142 355 148
rect 327 117 355 125
rect 372 139 389 170
rect 431 212 448 237
rect 431 162 448 170
rect 510 212 527 220
rect 510 162 527 170
rect 589 212 606 237
rect 589 162 606 170
rect 668 212 685 220
rect 668 162 685 170
rect 747 212 764 237
rect 747 162 764 170
rect 826 212 843 220
rect 775 141 809 149
rect 372 131 493 139
rect 389 114 465 131
rect 372 106 493 114
rect 248 91 276 99
rect 248 66 276 74
rect 327 91 355 99
rect 327 66 355 74
rect 214 -4 231 4
rect 293 46 310 54
rect 293 -21 310 4
rect 372 46 389 106
rect 589 69 628 86
rect 645 69 685 86
rect 589 54 685 69
rect 775 67 809 75
rect 905 212 922 237
rect 905 162 922 170
rect 984 212 1001 220
rect 984 162 1001 170
rect 1063 212 1080 237
rect 1063 162 1080 170
rect 372 -4 389 4
rect 431 46 448 54
rect 431 -21 448 4
rect 510 46 527 54
rect 510 -4 527 4
rect 589 46 606 54
rect 589 -4 606 4
rect 668 46 685 54
rect 668 -4 685 4
rect 747 46 764 54
rect 747 -4 764 4
rect 826 46 843 132
rect 826 -4 843 4
rect 905 69 944 86
rect 961 69 1001 86
rect 905 54 1001 69
rect 905 46 922 54
rect 905 -4 922 4
rect 984 46 1001 54
rect 984 -4 1001 4
rect 1063 46 1080 54
rect 1063 -4 1080 4
rect 589 -21 764 -4
rect 905 -21 1080 -4
rect -3 -43 1080 -38
rect -3 -60 9 -43
rect 1068 -60 1080 -43
<< viali >>
rect 214 243 1068 254
rect 1068 243 1080 254
rect 214 237 1080 243
rect 76 170 93 212
rect 36 123 54 140
rect -3 80 14 97
rect 115 80 133 97
rect 155 46 172 57
rect 155 40 172 46
rect 214 170 231 176
rect 214 159 231 170
rect 253 125 271 142
rect 332 148 350 165
rect 510 170 527 212
rect 668 170 685 212
rect 826 170 843 212
rect 372 114 389 131
rect 470 114 488 131
rect 253 74 271 91
rect 332 74 350 91
rect 772 75 775 109
rect 775 75 806 109
rect 826 132 843 170
rect 984 170 1001 212
rect 510 4 527 46
rect -3 -38 1080 -21
<< metal1 >>
rect 73 212 96 257
rect 185 254 1086 257
rect 185 237 214 254
rect 1080 237 1086 254
rect 185 234 1086 237
rect 510 215 527 218
rect 668 215 685 218
rect 73 170 76 212
rect 93 170 96 212
rect 507 212 530 215
rect 73 164 96 170
rect 211 176 356 182
rect 211 159 214 176
rect 231 165 356 176
rect 507 170 510 212
rect 527 170 530 212
rect 507 167 530 170
rect 665 212 688 215
rect 665 170 668 212
rect 685 170 688 212
rect 665 167 688 170
rect 823 212 846 218
rect 984 215 1001 218
rect 231 159 332 165
rect 211 153 234 159
rect 326 148 332 159
rect 350 148 356 165
rect 30 140 60 148
rect 326 145 356 148
rect 30 123 36 140
rect 54 123 60 140
rect 30 115 60 123
rect 247 142 312 145
rect 247 125 253 142
rect 271 131 312 142
rect 369 134 392 137
rect 369 131 494 134
rect 271 125 372 131
rect 247 122 372 125
rect 291 114 372 122
rect 389 114 470 131
rect 488 114 494 131
rect 369 111 494 114
rect 510 112 527 167
rect 668 112 685 167
rect 823 132 826 212
rect 843 166 846 212
rect 981 212 1004 215
rect 981 170 984 212
rect 1001 170 1004 212
rect 981 166 1004 170
rect 843 132 1119 166
rect 823 129 1119 132
rect 826 126 1119 129
rect 369 108 392 111
rect 510 109 1119 112
rect -6 100 17 103
rect -6 97 277 100
rect -6 80 -3 97
rect 14 80 115 97
rect 133 91 277 97
rect 133 80 253 91
rect -6 77 253 80
rect -6 74 17 77
rect 247 74 253 77
rect 271 74 277 91
rect 247 71 277 74
rect 326 91 356 94
rect 326 74 332 91
rect 350 74 356 91
rect 152 57 175 63
rect 326 57 356 74
rect 152 40 155 57
rect 172 40 356 57
rect 510 78 772 109
rect 510 72 628 78
rect 645 75 772 78
rect 806 75 1119 109
rect 645 72 1119 75
rect 510 49 527 72
rect 152 34 356 40
rect 507 46 530 49
rect 507 4 510 46
rect 527 4 530 46
rect 507 1 530 4
rect 510 -2 527 1
rect -9 -21 1086 -18
rect -9 -38 -3 -21
rect 1080 -38 1086 -21
rect -9 -41 1086 -38
<< labels >>
flabel metal1 30 115 60 148 0 FreeSans 160 0 0 0 in
port 1 nsew
flabel locali -3 122 14 139 0 FreeSans 80 90 0 0 in_b
flabel locali 155 116 172 143 0 FreeSans 80 90 0 0 in_bb
flabel locali 214 116 231 133 0 FreeSans 80 0 0 0 t2
flabel locali 372 80 389 97 0 FreeSans 80 0 0 0 t1
flabel metal1 1079 126 1119 166 0 FreeSans 160 0 0 0 out_b
port 2 nsew
flabel metal1 1079 72 1119 112 0 FreeSans 160 0 0 0 out
port 3 nsew
flabel metal1 73 234 96 257 0 FreeSans 160 0 0 0 vdd_l
port 4 nsew
flabel metal1 185 234 208 257 0 FreeSans 160 0 0 0 vdd_h
port 5 nsew
flabel metal1 -9 -41 14 -18 0 FreeSans 160 0 0 0 vss
port 6 nsew
<< end >>
