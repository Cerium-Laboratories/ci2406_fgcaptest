magic
tech sky130A
magscale 1 2
timestamp 1717172305
<< error_p >>
rect 80698 44914 81160 45074
rect 84698 44914 85160 45074
rect 88698 44914 89160 45074
rect 83064 44606 83528 44616
rect 87064 44606 87528 44616
rect 83064 44206 83528 44216
rect 87064 44206 87528 44216
rect 80698 43748 81160 43908
rect 84698 43748 85160 43908
rect 88698 43748 89160 43908
rect 80698 38914 81160 39074
rect 84698 38914 85160 39074
rect 88698 38914 89160 39074
rect 83064 38606 83528 38616
rect 87064 38606 87528 38616
rect 83064 38206 83528 38216
rect 87064 38206 87528 38216
rect 80698 37748 81160 37908
rect 84698 37748 85160 37908
rect 88698 37748 89160 37908
rect 80698 32914 81160 33074
rect 84698 32914 85160 33074
rect 88698 32914 89160 33074
rect 83064 32606 83528 32616
rect 87064 32606 87528 32616
rect 83064 32206 83528 32216
rect 87064 32206 87528 32216
rect 80698 31748 81160 31908
rect 84698 31748 85160 31908
rect 88698 31748 89160 31908
rect 80764 28748 81226 28908
rect 84764 28748 85226 28908
rect 88764 28748 89226 28908
rect 80764 10748 81226 10908
rect 84764 10748 85226 10908
rect 88764 10748 89226 10908
rect 92764 10748 93226 10908
rect 96764 10748 97226 10908
rect 100764 10748 101226 10908
rect 104764 10748 105226 10908
rect 108764 10748 109226 10908
rect 112764 10748 113226 10908
rect 116764 10748 117226 10908
rect 80764 7748 81226 7908
rect 84764 7748 85226 7908
rect 88764 7748 89226 7908
rect 92764 7748 93226 7908
rect 96764 7748 97226 7908
rect 100764 7748 101226 7908
rect 104764 7748 105226 7908
rect 108764 7748 109226 7908
rect 112764 7748 113226 7908
rect 116764 7748 117226 7908
rect 80764 4748 81226 4908
rect 84764 4748 85226 4908
rect 88764 4748 89226 4908
rect 92764 4748 93226 4908
rect 96764 4748 97226 4908
rect 100764 4748 101226 4908
rect 104764 4748 105226 4908
rect 108764 4748 109226 4908
rect 112764 4748 113226 4908
rect 116764 4748 117226 4908
rect 80764 1748 81226 1908
rect 84764 1748 85226 1908
rect 88764 1748 89226 1908
rect 92764 1748 93226 1908
rect 96764 1748 97226 1908
rect 100764 1748 101226 1908
rect 104764 1748 105226 1908
rect 108764 1748 109226 1908
rect 112764 1748 113226 1908
rect 116764 1748 117226 1908
<< error_s >>
rect 35319 -13380 35343 -13364
rect 35343 -13600 35346 -13380
rect 35651 -13742 35705 -13726
rect 35705 -13962 35708 -13742
rect 35961 -14056 36019 -14046
rect 36019 -14282 36028 -14056
rect 36291 -14382 36345 -14366
rect 51340 -14382 51345 -14366
rect 66340 -14382 66345 -14366
rect 36345 -14390 36348 -14382
rect 51345 -14390 51348 -14382
rect 66345 -14390 66348 -14382
rect 38597 -14642 38821 -14635
rect 53597 -14642 53821 -14635
rect 68597 -14642 68821 -14635
rect 38585 -14662 38597 -14642
rect 53585 -14662 53597 -14642
rect 68585 -14662 68597 -14642
rect 35085 -21555 35121 -21483
rect 35123 -21517 35157 -21483
rect 36614 -27109 36617 -27098
rect 51614 -27109 51617 -27098
rect 66614 -27109 66617 -27098
rect 36386 -27125 36614 -27109
rect 51386 -27125 51614 -27109
rect 66386 -27125 66614 -27109
rect 38854 -27378 38857 -27158
rect 53854 -27378 53857 -27158
rect 68854 -27378 68857 -27158
rect 36291 -27432 36294 -27380
rect 38857 -27394 38860 -27378
rect 53857 -27394 53860 -27378
rect 68857 -27394 68860 -27378
rect 36058 -27448 36291 -27432
rect 35971 -27752 35974 -27698
rect 35854 -27768 35971 -27752
rect 35651 -28072 35654 -28018
rect 35418 -28088 35651 -28072
rect 35319 -28396 35332 -28380
use array_core  array_core_0
timestamp 1717172305
transform 1 0 40000 0 1 0
box -40000 0 80032 89628
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1716601000
transform -1 0 37600 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_2
timestamp 1716601000
transform -1 0 67600 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_3
timestamp 1716601000
transform -1 0 52600 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__analog_minesd_pad_short  sky130_ef_io__analog_minesd_pad_short_4
timestamp 1716601000
transform -1 0 82600 0 -1 6200
box 0 14007 15000 40000
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1716601000
transform 1 0 8540 0 1 -25060
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_1
timestamp 1716601000
transform 1 0 106540 0 1 -23060
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_2
timestamp 1716601000
transform 1 0 84540 0 1 -21660
box -540 -540 12540 14540
<< end >>
