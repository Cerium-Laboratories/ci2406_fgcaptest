magic
tech sky130A
timestamp 1716945357
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vin
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 vout
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 en
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 en_b
port 3 nsew
<< end >>
