** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/test_diffamp_nmos.sch
**.subckt test_diffamp_nmos
VDD VDD GND {VDD}
vb vb GND {VBIAS}
v1 v1 GND 3 pwl(0 3 1u 3 1.1u 4.7 1.5u 4 1.7u 0.5 2u 0.1 2.1u 3)
v2 v2 GND 2
R1 vout GND 1T m=1
x1 v1 vout vb vout VDD GND diffamp_nmos
C1 vout GND 26f m=1
**** begin user architecture code
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.options reltol=0.0001 abstol=10e-15
.include diffamp_nmos.spice
.param VDD=5
.param VSS=0
.param VBIAS=1
.options savecurrents
* .options reltol=0.01 abstol=10e-12
.control
  save all
  op
  remzerovec
  write test_diffamp_nmos.raw
  set appendwrite
  * vb sweep
  dc v1 0 6 0.2 vb 0 5 1
  remzerovec
  write test_diffamp_nmos.raw
  * dc sweep
  dc v1 0 5 0.1
  remzerovec
  write test_diffamp_nmos.raw
  * tran
  tran 1n 3u
  remzerovec
  write test_diffamp_nmos.raw
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
