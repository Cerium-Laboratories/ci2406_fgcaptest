magic
tech sky130A
timestamp 1717695944
<< metal1 >>
rect 32441 1980 32519 1983
rect 25998 1977 32441 1980
rect 25998 1951 26014 1977
rect 26066 1951 26814 1977
rect 26866 1951 27614 1977
rect 27666 1951 28414 1977
rect 28466 1951 29214 1977
rect 29266 1951 30014 1977
rect 30066 1951 30814 1977
rect 30866 1951 31614 1977
rect 31666 1951 32441 1977
rect 25998 1900 32441 1951
rect 26180 1854 26238 1857
rect 26180 1802 26183 1854
rect 26235 1802 26238 1854
rect 26373 1844 26415 1900
rect 26580 1854 26638 1857
rect 26180 1799 26238 1802
rect 26580 1802 26583 1854
rect 26635 1802 26638 1854
rect 26773 1844 26815 1900
rect 26980 1854 27038 1857
rect 26580 1799 26638 1802
rect 26980 1802 26983 1854
rect 27035 1802 27038 1854
rect 27173 1844 27215 1900
rect 27380 1854 27438 1857
rect 26980 1799 27038 1802
rect 27380 1802 27383 1854
rect 27435 1802 27438 1854
rect 27573 1844 27615 1900
rect 27780 1854 27838 1857
rect 27380 1799 27438 1802
rect 27780 1802 27783 1854
rect 27835 1802 27838 1854
rect 27973 1844 28015 1900
rect 28180 1854 28238 1857
rect 27780 1799 27838 1802
rect 28180 1802 28183 1854
rect 28235 1802 28238 1854
rect 28373 1844 28415 1900
rect 28580 1854 28638 1857
rect 28180 1799 28238 1802
rect 28580 1802 28583 1854
rect 28635 1802 28638 1854
rect 28773 1844 28815 1900
rect 28980 1854 29038 1857
rect 28580 1799 28638 1802
rect 28980 1802 28983 1854
rect 29035 1802 29038 1854
rect 29173 1844 29215 1900
rect 29380 1854 29438 1857
rect 28980 1799 29038 1802
rect 29380 1802 29383 1854
rect 29435 1802 29438 1854
rect 29573 1844 29615 1900
rect 29780 1854 29838 1857
rect 29380 1799 29438 1802
rect 29780 1802 29783 1854
rect 29835 1802 29838 1854
rect 29973 1844 30015 1900
rect 30180 1854 30238 1857
rect 29780 1799 29838 1802
rect 30180 1802 30183 1854
rect 30235 1802 30238 1854
rect 30373 1844 30415 1900
rect 30580 1854 30638 1857
rect 30180 1799 30238 1802
rect 30580 1802 30583 1854
rect 30635 1802 30638 1854
rect 30773 1844 30815 1900
rect 30980 1854 31038 1857
rect 30580 1799 30638 1802
rect 30980 1802 30983 1854
rect 31035 1802 31038 1854
rect 31173 1844 31215 1900
rect 31380 1854 31438 1857
rect 30980 1799 31038 1802
rect 31380 1802 31383 1854
rect 31435 1802 31438 1854
rect 31573 1844 31615 1900
rect 31780 1854 31838 1857
rect 31380 1799 31438 1802
rect 31780 1802 31783 1854
rect 31835 1802 31838 1854
rect 31973 1844 32015 1900
rect 32180 1854 32238 1857
rect 31780 1799 31838 1802
rect 32180 1802 32183 1854
rect 32235 1802 32238 1854
rect 32373 1844 32415 1900
rect 32441 1897 32519 1900
rect 32180 1799 32238 1802
rect 53000 -10220 53130 -10200
rect 53000 -13890 53010 -10220
rect 53110 -13890 53130 -10220
rect 53000 -13910 53130 -13890
<< via1 >>
rect 26014 2130 26066 2156
rect 26814 2130 26866 2156
rect 27614 2130 27666 2156
rect 28414 2130 28466 2156
rect 29214 2130 29266 2156
rect 30014 2130 30066 2156
rect 30814 2130 30866 2156
rect 31614 2130 31666 2156
rect 26014 1951 26066 1977
rect 26814 1951 26866 1977
rect 27614 1951 27666 1977
rect 28414 1951 28466 1977
rect 29214 1951 29266 1977
rect 30014 1951 30066 1977
rect 30814 1951 30866 1977
rect 31614 1951 31666 1977
rect 32441 1900 32519 1980
rect 26183 1802 26235 1854
rect 26583 1802 26635 1854
rect 26983 1802 27035 1854
rect 27383 1802 27435 1854
rect 27783 1802 27835 1854
rect 28183 1802 28235 1854
rect 28583 1802 28635 1854
rect 28983 1802 29035 1854
rect 29383 1802 29435 1854
rect 29783 1802 29835 1854
rect 30183 1802 30235 1854
rect 30583 1802 30635 1854
rect 30983 1802 31035 1854
rect 31383 1802 31435 1854
rect 31783 1802 31835 1854
rect 32183 1802 32235 1854
rect 53010 -13890 53110 -10220
<< metal2 >>
rect 26011 2156 26069 2159
rect 26011 2130 26014 2156
rect 26066 2130 26069 2156
rect 26011 1977 26069 2130
rect 26811 2156 26869 2159
rect 26811 2130 26814 2156
rect 26866 2130 26869 2156
rect 26011 1951 26014 1977
rect 26066 1951 26069 1977
rect 26011 1948 26069 1951
rect 26180 1854 26238 2000
rect 26180 1802 26183 1854
rect 26235 1802 26238 1854
rect 26180 1799 26238 1802
rect 26580 1854 26638 2000
rect 26811 1977 26869 2130
rect 27611 2156 27669 2159
rect 27611 2130 27614 2156
rect 27666 2130 27669 2156
rect 26811 1951 26814 1977
rect 26866 1951 26869 1977
rect 26811 1948 26869 1951
rect 26580 1802 26583 1854
rect 26635 1802 26638 1854
rect 26580 1799 26638 1802
rect 26980 1854 27038 2000
rect 26980 1802 26983 1854
rect 27035 1802 27038 1854
rect 26980 1799 27038 1802
rect 27380 1854 27438 2000
rect 27611 1977 27669 2130
rect 28411 2156 28469 2159
rect 28411 2130 28414 2156
rect 28466 2130 28469 2156
rect 27611 1951 27614 1977
rect 27666 1951 27669 1977
rect 27611 1948 27669 1951
rect 27380 1802 27383 1854
rect 27435 1802 27438 1854
rect 27380 1799 27438 1802
rect 27780 1854 27838 2000
rect 27780 1802 27783 1854
rect 27835 1802 27838 1854
rect 27780 1799 27838 1802
rect 28180 1854 28238 2000
rect 28411 1977 28469 2130
rect 29211 2156 29269 2159
rect 29211 2130 29214 2156
rect 29266 2130 29269 2156
rect 28411 1951 28414 1977
rect 28466 1951 28469 1977
rect 28411 1948 28469 1951
rect 28180 1802 28183 1854
rect 28235 1802 28238 1854
rect 28180 1799 28238 1802
rect 28580 1854 28638 2000
rect 28580 1802 28583 1854
rect 28635 1802 28638 1854
rect 28580 1799 28638 1802
rect 28980 1854 29038 2000
rect 29211 1977 29269 2130
rect 30011 2156 30069 2159
rect 30011 2130 30014 2156
rect 30066 2130 30069 2156
rect 29211 1951 29214 1977
rect 29266 1951 29269 1977
rect 29211 1948 29269 1951
rect 28980 1802 28983 1854
rect 29035 1802 29038 1854
rect 28980 1799 29038 1802
rect 29380 1854 29438 2000
rect 29380 1802 29383 1854
rect 29435 1802 29438 1854
rect 29380 1799 29438 1802
rect 29780 1854 29838 2000
rect 30011 1977 30069 2130
rect 30811 2156 30869 2159
rect 30811 2130 30814 2156
rect 30866 2130 30869 2156
rect 30011 1951 30014 1977
rect 30066 1951 30069 1977
rect 30011 1948 30069 1951
rect 29780 1802 29783 1854
rect 29835 1802 29838 1854
rect 29780 1799 29838 1802
rect 30180 1854 30238 2000
rect 30180 1802 30183 1854
rect 30235 1802 30238 1854
rect 30180 1799 30238 1802
rect 30580 1854 30638 2000
rect 30811 1977 30869 2130
rect 31611 2156 31669 2159
rect 31611 2130 31614 2156
rect 31666 2130 31669 2156
rect 30811 1951 30814 1977
rect 30866 1951 30869 1977
rect 30811 1948 30869 1951
rect 30580 1802 30583 1854
rect 30635 1802 30638 1854
rect 30580 1799 30638 1802
rect 30980 1854 31038 2000
rect 30980 1802 30983 1854
rect 31035 1802 31038 1854
rect 30980 1799 31038 1802
rect 31380 1854 31438 2000
rect 31611 1977 31669 2130
rect 31611 1951 31614 1977
rect 31666 1951 31669 1977
rect 31611 1948 31669 1951
rect 31380 1802 31383 1854
rect 31435 1802 31438 1854
rect 31380 1799 31438 1802
rect 31780 1854 31838 2000
rect 31780 1802 31783 1854
rect 31835 1802 31838 1854
rect 31780 1799 31838 1802
rect 32180 1854 32238 2000
rect 32441 1980 32519 2130
rect 32441 1897 32519 1900
rect 32180 1802 32183 1854
rect 32235 1802 32238 1854
rect 32180 1799 32238 1802
rect 53000 -10220 53130 -10200
rect 53000 -13890 53010 -10220
rect 53110 -13890 53130 -10220
rect 53000 -13910 53130 -13890
<< via2 >>
rect 53010 -13890 53110 -10220
<< metal3 >>
rect 27300 45500 27500 45600
rect 27900 45500 28100 45600
rect 28500 45500 28700 45600
rect 29100 45500 29300 45600
rect 29700 45500 29900 45600
rect 30300 45500 30500 45600
rect 30900 45500 31100 45600
rect 31500 45500 31700 45600
rect 32100 45500 32300 45600
rect 7200 -2410 22750 -2400
rect 7200 -2990 7210 -2410
rect 7790 -2990 22750 -2410
rect 7200 -3000 22750 -2990
rect 22860 -3100 23520 -2600
rect 14700 -3110 23520 -3100
rect 14700 -3690 14710 -3110
rect 15290 -3690 23520 -3110
rect 14700 -3700 23520 -3690
rect 24400 -3900 24800 -2600
rect 22200 -3910 24800 -3900
rect 22200 -4290 22210 -3910
rect 22790 -4290 24800 -3910
rect 22200 -4300 24800 -4290
rect 37200 -3910 37800 -2600
rect 43900 -2620 46100 -2600
rect 43900 -2880 43920 -2620
rect 46080 -2880 46100 -2620
rect 43900 -2900 46100 -2880
rect 37200 -4290 37210 -3910
rect 37790 -4290 37800 -3910
rect 37200 -4310 37800 -4290
rect 47960 -10220 53130 -10200
rect 47960 -13890 53010 -10220
rect 53110 -13890 53130 -10220
rect 47960 -13910 53130 -13890
<< via3 >>
rect 7210 -2990 7790 -2410
rect 14710 -3690 15290 -3110
rect 22210 -4290 22790 -3910
rect 43920 -2880 46080 -2620
rect 37210 -4290 37790 -3910
<< metal4 >>
rect -4800 45200 24900 45600
rect -4800 -17400 -4400 45200
rect 24100 43900 24900 45200
rect 60060 43680 63300 43700
rect 60060 43320 60080 43680
rect 60440 43320 63300 43680
rect 60060 43300 63300 43320
rect 62900 33700 63300 43300
rect 60060 33680 63300 33700
rect 60060 33320 60080 33680
rect 60440 33320 63300 33680
rect 60060 33300 63300 33320
rect 62900 23700 63300 33300
rect 60060 23680 63300 23700
rect 60060 23320 60080 23680
rect 60440 23320 63300 23680
rect 60060 23300 63300 23320
rect 62900 13700 63300 23300
rect 60060 13680 63300 13700
rect 60060 13320 60080 13680
rect 60440 13320 63300 13680
rect 60060 13300 63300 13320
rect 62900 3700 63300 13300
rect 60060 3680 63300 3700
rect 60060 3320 60080 3680
rect 60440 3320 63300 3680
rect 60060 3300 63300 3320
rect 7000 -2410 8000 -2400
rect 7000 -2990 7210 -2410
rect 7790 -2990 8000 -2410
rect 7000 -6600 8000 -2990
rect 14500 -3110 15500 -3100
rect 14500 -3690 14710 -3110
rect 15290 -3690 15500 -3110
rect 14500 -6600 15500 -3690
rect 22000 -3910 23000 -3900
rect 22000 -4290 22210 -3910
rect 22790 -4290 23000 -3910
rect 22000 -6700 23000 -4290
rect 29000 -4500 31000 -2600
rect 43900 -2620 46100 -2600
rect 43900 -2880 43920 -2620
rect 46080 -2880 46100 -2620
rect 43900 -2900 46100 -2880
rect 37000 -3910 38000 -3900
rect 37000 -4290 37210 -3910
rect 37790 -4290 38000 -3910
rect 29080 -6900 30939 -4500
rect 37000 -6700 38000 -4290
rect 62900 -6300 63300 3300
rect 60060 -6320 63300 -6300
rect 60060 -6680 60080 -6320
rect 60440 -6680 63300 -6320
rect 60060 -6700 63300 -6680
rect 62900 -17000 63300 -6700
rect 60060 -17020 63300 -17000
rect 60060 -17380 60080 -17020
rect 60440 -17380 63300 -17020
rect 60060 -17400 63300 -17380
<< via4 >>
rect 60080 43320 60440 43680
rect 60080 33320 60440 33680
rect 60080 23320 60440 23680
rect 60080 13320 60440 13680
rect 60080 3320 60440 3680
rect 43920 -2880 46080 -2620
rect 60080 -6680 60440 -6320
rect 60080 -17380 60440 -17020
<< metal5 >>
rect -500 43300 -100 43700
rect 60060 43680 60460 43700
rect 60060 43320 60080 43680
rect 60440 43320 60460 43680
rect 60060 43300 60460 43320
rect 60060 33680 60460 33700
rect 60060 33320 60080 33680
rect 60440 33320 60460 33680
rect 60060 33300 60460 33320
rect 60060 23680 60460 23700
rect 60060 23320 60080 23680
rect 60440 23320 60460 23680
rect 60060 23300 60460 23320
rect 60060 13680 60460 13700
rect 60060 13320 60080 13680
rect 60440 13320 60460 13680
rect 60060 13300 60460 13320
rect 60060 3680 60460 3700
rect 60060 3320 60080 3680
rect 60440 3320 60460 3680
rect 60060 3300 60460 3320
rect -500 -15400 -100 -1500
rect 43900 -2620 46100 -2600
rect 43900 -2880 43920 -2620
rect 46080 -2880 46100 -2620
rect 43900 -7300 46100 -2880
rect 54400 -7010 56600 -2600
rect 60060 -6320 60460 -1000
rect 60060 -6680 60080 -6320
rect 60440 -6680 60460 -6320
rect 4755 -14198 10250 -7687
rect 12255 -14198 17750 -7687
rect 19755 -14198 25250 -7687
rect 27255 -14198 32750 -7687
rect 34755 -14198 40250 -7687
rect 41860 -14580 48140 -7300
rect 52360 -14580 58640 -7300
rect 41730 -14980 48270 -14710
rect 41250 -15400 48270 -14980
rect 60060 -15400 60460 -6680
rect -500 -17020 60460 -15400
rect -500 -17380 60080 -17020
rect 60440 -17380 60460 -17020
rect -500 -17400 60460 -17380
use array_core  array_core_0
timestamp 1717695944
transform 1 0 20000 0 1 0
box -20500 -2600 40460 45600
use bare_pad_gnd  bare_pad_gnd_0
timestamp 1717628967
transform 1 0 41730 0 1 -14710
box 0 0 6540 7540
use vtun_pad  vtun_pad_0
timestamp 1717630197
transform 1 0 34200 0 1 -14700
box 0 0 6540 8100
use vtun_pad  vtun_pad_1
timestamp 1717630197
transform 1 0 52230 0 1 -14710
box 0 0 6540 8100
use vtun_pad  vtun_pad_2
timestamp 1717630197
transform 1 0 4200 0 1 -14700
box 0 0 6540 8100
use vtun_pad  vtun_pad_3
timestamp 1717630197
transform 1 0 11700 0 1 -14700
box 0 0 6540 8100
use vtun_pad  vtun_pad_4
timestamp 1717630197
transform 1 0 19200 0 1 -14700
box 0 0 6540 8100
use vtun_pad  vtun_pad_5
timestamp 1717630197
transform 1 0 26700 0 1 -14700
box 0 0 6540 8100
<< labels >>
flabel metal5 41860 -14580 48140 -7300 0 FreeSans 3200 0 0 0 VGND
flabel metal5 19755 -14198 25250 -7687 0 FreeSans 3200 0 0 0 VOUT0
flabel metal5 34755 -14198 40250 -7687 0 FreeSans 3200 0 0 0 VOUT1
flabel metal5 27255 -14198 32750 -7687 0 FreeSans 3200 0 0 0 VINJ
flabel metal5 12255 -14198 17750 -7687 0 FreeSans 3200 0 0 0 VCTRL
flabel metal5 4755 -14198 10250 -7687 0 FreeSans 3200 0 0 0 VSRC
flabel metal5 52360 -14580 58640 -7300 0 FreeSans 3200 0 0 0 VTUN
flabel metal3 27300 45500 27500 45600 0 FreeSans 400 0 0 0 addr[0]
port 3 n signal input
flabel metal3 27900 45500 28100 45600 0 FreeSans 400 0 0 0 addr[1]
port 4 n signal input
flabel metal3 28500 45500 28700 45600 0 FreeSans 400 0 0 0 addr[2]
port 5 n signal input
flabel metal3 29100 45500 29300 45600 0 FreeSans 400 0 0 0 addr[3]
port 6 n signal input
flabel metal3 29700 45500 29900 45600 0 FreeSans 400 0 0 0 addr[4]
port 7 n signal input
flabel metal3 30300 45500 30500 45600 0 FreeSans 400 0 0 0 addr[5]
port 8 n signal input
flabel metal3 30900 45500 31100 45600 0 FreeSans 400 0 0 0 addr[6]
port 9 n signal input
flabel metal3 31500 45500 31700 45600 0 FreeSans 400 0 0 0 addr[7]
port 10 n signal input
flabel metal3 32100 45500 32300 45600 0 FreeSans 400 0 0 0 addr[8]
port 11 n signal input
flabel metal4 62900 -17400 63300 43700 0 FreeSans 1600 180 0 0 vssd2
port 13 nsew ground bidirectional abutment
flabel metal4 -4800 -6800 -4400 45600 0 FreeSans 1600 0 0 0 vccd2
port 14 nsew power bidirectional abutment
<< properties >>
string FIXE_BBOX -9600 -34800 126600 91200 
string FIXED_BBOX -4800 -17400 63300 45600
<< end >>
