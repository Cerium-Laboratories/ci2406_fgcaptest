magic
tech sky130A
timestamp 1717011964
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vinj
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 vinj_en_b
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 vtun
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 vctrl
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 vsrc
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 VGND
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 vfg
port 6 nsew
<< end >>
