magic
tech sky130A
timestamp 1717172305
<< error_p >>
rect 20382 5374 20613 5454
rect 22382 5374 22613 5454
rect 24382 5374 24613 5454
rect 26382 5374 26613 5454
rect 28382 5374 28613 5454
rect 30382 5374 30613 5454
rect 32382 5374 32613 5454
rect 34382 5374 34613 5454
rect 36382 5374 36613 5454
rect 38382 5374 38613 5454
rect 20382 3874 20613 3954
rect 22382 3874 22613 3954
rect 24382 3874 24613 3954
rect 26382 3874 26613 3954
rect 28382 3874 28613 3954
rect 30382 3874 30613 3954
rect 32382 3874 32613 3954
rect 34382 3874 34613 3954
rect 36382 3874 36613 3954
rect 38382 3874 38613 3954
rect 20382 2374 20613 2454
rect 22382 2374 22613 2454
rect 24382 2374 24613 2454
rect 26382 2374 26613 2454
rect 28382 2374 28613 2454
rect 30382 2374 30613 2454
rect 32382 2374 32613 2454
rect 34382 2374 34613 2454
rect 36382 2374 36613 2454
rect 38382 2374 38613 2454
rect 20382 874 20613 954
rect 22382 874 22613 954
rect 24382 874 24613 954
rect 26382 874 26613 954
rect 28382 874 28613 954
rect 30382 874 30613 954
rect 32382 874 32613 954
rect 34382 874 34613 954
rect 36382 874 36613 954
rect 38382 874 38613 954
<< error_s >>
rect 20349 22457 20580 22537
rect 22349 22457 22580 22537
rect 24349 22457 24580 22537
rect 21532 22303 21764 22308
rect 23532 22303 23764 22308
rect 21532 22103 21764 22108
rect 23532 22103 23764 22108
rect 20349 21874 20580 21954
rect 22349 21874 22580 21954
rect 24349 21874 24580 21954
rect 20349 19457 20580 19537
rect 22349 19457 22580 19537
rect 24349 19457 24580 19537
rect 21532 19303 21764 19308
rect 23532 19303 23764 19308
rect 21532 19103 21764 19108
rect 23532 19103 23764 19108
rect 20349 18874 20580 18954
rect 22349 18874 22580 18954
rect 24349 18874 24580 18954
rect 20349 16457 20580 16537
rect 22349 16457 22580 16537
rect 24349 16457 24580 16537
rect 21532 16303 21764 16308
rect 23532 16303 23764 16308
rect 21532 16103 21764 16108
rect 23532 16103 23764 16108
rect 20349 15874 20580 15954
rect 22349 15874 22580 15954
rect 24349 15874 24580 15954
rect 20382 14374 20613 14454
rect 22382 14374 22613 14454
rect 24382 14374 24613 14454
<< metal1 >>
rect 4897 41793 4900 41871
rect 4980 41793 4983 41871
rect 14597 41793 14600 41871
rect 14680 41793 14683 41871
rect 4900 41767 4980 41793
rect 4844 41725 4980 41767
rect 4799 41587 4857 41590
rect 4799 41535 4802 41587
rect 4854 41535 4857 41587
rect 4799 41532 4857 41535
rect 4900 41367 4980 41725
rect 4844 41325 4980 41367
rect 4799 41187 4857 41190
rect 4799 41135 4802 41187
rect 4854 41135 4857 41187
rect 4799 41132 4857 41135
rect 4900 41018 4980 41325
rect 14600 41767 14680 41793
rect 14600 41725 14736 41767
rect 14600 41367 14680 41725
rect 14723 41587 14781 41590
rect 14723 41535 14726 41587
rect 14778 41535 14781 41587
rect 14723 41532 14781 41535
rect 14600 41325 14736 41367
rect 14600 41018 14680 41325
rect 14723 41187 14781 41190
rect 14723 41135 14726 41187
rect 14778 41135 14781 41187
rect 14723 41132 14781 41135
rect 4900 40967 4951 41018
rect 4844 40966 4951 40967
rect 4977 40966 4980 41018
rect 14600 40966 14603 41018
rect 14629 40967 14680 41018
rect 14629 40966 14736 40967
rect 4844 40925 4980 40966
rect 4799 40787 4857 40790
rect 4799 40735 4802 40787
rect 4854 40735 4857 40787
rect 4799 40732 4857 40735
rect 4900 40567 4980 40925
rect 4844 40525 4980 40567
rect 4799 40387 4857 40390
rect 4799 40335 4802 40387
rect 4854 40335 4857 40387
rect 4799 40332 4857 40335
rect 4900 40218 4980 40525
rect 14600 40925 14736 40966
rect 14600 40567 14680 40925
rect 14723 40787 14781 40790
rect 14723 40735 14726 40787
rect 14778 40735 14781 40787
rect 14723 40732 14781 40735
rect 14600 40525 14736 40567
rect 14600 40218 14680 40525
rect 14723 40387 14781 40390
rect 14723 40335 14726 40387
rect 14778 40335 14781 40387
rect 14723 40332 14781 40335
rect 4900 40167 4951 40218
rect 4844 40166 4951 40167
rect 4977 40166 4980 40218
rect 14600 40166 14603 40218
rect 14629 40167 14680 40218
rect 14629 40166 14736 40167
rect 4844 40125 4980 40166
rect 4799 39987 4857 39990
rect 4799 39935 4802 39987
rect 4854 39935 4857 39987
rect 4799 39932 4857 39935
rect 4900 39767 4980 40125
rect 4844 39725 4980 39767
rect 4799 39587 4857 39590
rect 4799 39535 4802 39587
rect 4854 39535 4857 39587
rect 4799 39532 4857 39535
rect 4900 39418 4980 39725
rect 14600 40125 14736 40166
rect 14600 39767 14680 40125
rect 14723 39987 14781 39990
rect 14723 39935 14726 39987
rect 14778 39935 14781 39987
rect 14723 39932 14781 39935
rect 14600 39725 14736 39767
rect 14600 39418 14680 39725
rect 14723 39587 14781 39590
rect 14723 39535 14726 39587
rect 14778 39535 14781 39587
rect 14723 39532 14781 39535
rect 4900 39367 4951 39418
rect 4844 39366 4951 39367
rect 4977 39366 4980 39418
rect 14600 39366 14603 39418
rect 14629 39367 14680 39418
rect 14629 39366 14736 39367
rect 4844 39325 4980 39366
rect 4799 39187 4857 39190
rect 4799 39135 4802 39187
rect 4854 39135 4857 39187
rect 4799 39132 4857 39135
rect 4900 38967 4980 39325
rect 4844 38925 4980 38967
rect 4799 38787 4857 38790
rect 4799 38735 4802 38787
rect 4854 38735 4857 38787
rect 4799 38732 4857 38735
rect 4900 38618 4980 38925
rect 14600 39325 14736 39366
rect 14600 38967 14680 39325
rect 14723 39187 14781 39190
rect 14723 39135 14726 39187
rect 14778 39135 14781 39187
rect 14723 39132 14781 39135
rect 14600 38925 14736 38967
rect 14600 38618 14680 38925
rect 14723 38787 14781 38790
rect 14723 38735 14726 38787
rect 14778 38735 14781 38787
rect 14723 38732 14781 38735
rect 4900 38567 4951 38618
rect 4844 38566 4951 38567
rect 4977 38566 4980 38618
rect 14600 38566 14603 38618
rect 14629 38567 14680 38618
rect 14629 38566 14736 38567
rect 4844 38525 4980 38566
rect 4799 38387 4857 38390
rect 4799 38335 4802 38387
rect 4854 38335 4857 38387
rect 4799 38332 4857 38335
rect 4900 38167 4980 38525
rect 4844 38125 4980 38167
rect 4799 37987 4857 37990
rect 4799 37935 4802 37987
rect 4854 37935 4857 37987
rect 4799 37932 4857 37935
rect 4900 37818 4980 38125
rect 14600 38525 14736 38566
rect 14600 38167 14680 38525
rect 14723 38387 14781 38390
rect 14723 38335 14726 38387
rect 14778 38335 14781 38387
rect 14723 38332 14781 38335
rect 14600 38125 14736 38167
rect 14600 37818 14680 38125
rect 14723 37987 14781 37990
rect 14723 37935 14726 37987
rect 14778 37935 14781 37987
rect 14723 37932 14781 37935
rect 4900 37767 4951 37818
rect 4844 37766 4951 37767
rect 4977 37766 4980 37818
rect 14600 37766 14603 37818
rect 14629 37767 14680 37818
rect 14629 37766 14736 37767
rect 4844 37725 4980 37766
rect 4799 37587 4857 37590
rect 4799 37535 4802 37587
rect 4854 37535 4857 37587
rect 4799 37532 4857 37535
rect 4900 37367 4980 37725
rect 4844 37325 4980 37367
rect 4799 37187 4857 37190
rect 4799 37135 4802 37187
rect 4854 37135 4857 37187
rect 4799 37132 4857 37135
rect 4900 37018 4980 37325
rect 14600 37725 14736 37766
rect 14600 37367 14680 37725
rect 14723 37587 14781 37590
rect 14723 37535 14726 37587
rect 14778 37535 14781 37587
rect 14723 37532 14781 37535
rect 14600 37325 14736 37367
rect 14600 37018 14680 37325
rect 14723 37187 14781 37190
rect 14723 37135 14726 37187
rect 14778 37135 14781 37187
rect 14723 37132 14781 37135
rect 4900 36967 4951 37018
rect 4844 36966 4951 36967
rect 4977 36966 4980 37018
rect 14600 36966 14603 37018
rect 14629 36967 14680 37018
rect 14629 36966 14736 36967
rect 4844 36925 4980 36966
rect 4799 36787 4857 36790
rect 4799 36735 4802 36787
rect 4854 36735 4857 36787
rect 4799 36732 4857 36735
rect 4900 36567 4980 36925
rect 4844 36525 4980 36567
rect 4799 36387 4857 36390
rect 4799 36335 4802 36387
rect 4854 36335 4857 36387
rect 4799 36332 4857 36335
rect 4900 36218 4980 36525
rect 14600 36925 14736 36966
rect 14600 36567 14680 36925
rect 14723 36787 14781 36790
rect 14723 36735 14726 36787
rect 14778 36735 14781 36787
rect 14723 36732 14781 36735
rect 14600 36525 14736 36567
rect 14600 36218 14680 36525
rect 14723 36387 14781 36390
rect 14723 36335 14726 36387
rect 14778 36335 14781 36387
rect 14723 36332 14781 36335
rect 4900 36167 4951 36218
rect 4844 36166 4951 36167
rect 4977 36166 4980 36218
rect 14600 36166 14603 36218
rect 14629 36167 14680 36218
rect 14629 36166 14736 36167
rect 4844 36125 4980 36166
rect 4799 35987 4857 35990
rect 4799 35935 4802 35987
rect 4854 35935 4857 35987
rect 4799 35932 4857 35935
rect 4900 35767 4980 36125
rect 4844 35725 4980 35767
rect 4799 35587 4857 35590
rect 4799 35535 4802 35587
rect 4854 35535 4857 35587
rect 4799 35532 4857 35535
rect 4900 35418 4980 35725
rect 14600 36125 14736 36166
rect 14600 35767 14680 36125
rect 14723 35987 14781 35990
rect 14723 35935 14726 35987
rect 14778 35935 14781 35987
rect 14723 35932 14781 35935
rect 14600 35725 14736 35767
rect 14600 35418 14680 35725
rect 14723 35587 14781 35590
rect 14723 35535 14726 35587
rect 14778 35535 14781 35587
rect 14723 35532 14781 35535
rect 4900 35367 4951 35418
rect 4844 35366 4951 35367
rect 4977 35366 4980 35418
rect 14600 35366 14603 35418
rect 14629 35367 14680 35418
rect 14629 35366 14736 35367
rect 4844 35325 4980 35366
rect 4799 35187 4857 35190
rect 4799 35135 4802 35187
rect 4854 35135 4857 35187
rect 4799 35132 4857 35135
rect 4900 34967 4980 35325
rect 4844 34925 4980 34967
rect 4799 34787 4857 34790
rect 4799 34735 4802 34787
rect 4854 34735 4857 34787
rect 4799 34732 4857 34735
rect 4900 34618 4980 34925
rect 14600 35325 14736 35366
rect 14600 34967 14680 35325
rect 14723 35187 14781 35190
rect 14723 35135 14726 35187
rect 14778 35135 14781 35187
rect 14723 35132 14781 35135
rect 14600 34925 14736 34967
rect 14600 34618 14680 34925
rect 14723 34787 14781 34790
rect 14723 34735 14726 34787
rect 14778 34735 14781 34787
rect 14723 34732 14781 34735
rect 4900 34567 4951 34618
rect 4844 34566 4951 34567
rect 4977 34566 4980 34618
rect 14600 34566 14603 34618
rect 14629 34567 14680 34618
rect 14629 34566 14736 34567
rect 4844 34525 4980 34566
rect 4799 34387 4857 34390
rect 4799 34335 4802 34387
rect 4854 34335 4857 34387
rect 4799 34332 4857 34335
rect 4900 34167 4980 34525
rect 4844 34125 4980 34167
rect 4799 33987 4857 33990
rect 4799 33935 4802 33987
rect 4854 33935 4857 33987
rect 4799 33932 4857 33935
rect 4900 33818 4980 34125
rect 14600 34525 14736 34566
rect 14600 34167 14680 34525
rect 14723 34387 14781 34390
rect 14723 34335 14726 34387
rect 14778 34335 14781 34387
rect 14723 34332 14781 34335
rect 14600 34125 14736 34167
rect 14600 33818 14680 34125
rect 14723 33987 14781 33990
rect 14723 33935 14726 33987
rect 14778 33935 14781 33987
rect 14723 33932 14781 33935
rect 4900 33767 4951 33818
rect 4844 33766 4951 33767
rect 4977 33766 4980 33818
rect 14600 33766 14603 33818
rect 14629 33767 14680 33818
rect 14629 33766 14736 33767
rect 4844 33725 4980 33766
rect 4799 33587 4857 33590
rect 4799 33535 4802 33587
rect 4854 33535 4857 33587
rect 4799 33532 4857 33535
rect 4900 33367 4980 33725
rect 4844 33325 4980 33367
rect 4799 33187 4857 33190
rect 4799 33135 4802 33187
rect 4854 33135 4857 33187
rect 4799 33132 4857 33135
rect 4900 33018 4980 33325
rect 14600 33725 14736 33766
rect 14600 33367 14680 33725
rect 14723 33587 14781 33590
rect 14723 33535 14726 33587
rect 14778 33535 14781 33587
rect 14723 33532 14781 33535
rect 14600 33325 14736 33367
rect 14600 33018 14680 33325
rect 14723 33187 14781 33190
rect 14723 33135 14726 33187
rect 14778 33135 14781 33187
rect 14723 33132 14781 33135
rect 4900 32967 4951 33018
rect 4844 32966 4951 32967
rect 4977 32966 4980 33018
rect 14600 32966 14603 33018
rect 14629 32967 14680 33018
rect 14629 32966 14736 32967
rect 4844 32925 4980 32966
rect 4799 32787 4857 32790
rect 4799 32735 4802 32787
rect 4854 32735 4857 32787
rect 4799 32732 4857 32735
rect 4900 32567 4980 32925
rect 4844 32525 4980 32567
rect 4799 32387 4857 32390
rect 4799 32335 4802 32387
rect 4854 32335 4857 32387
rect 4799 32332 4857 32335
rect 4900 32218 4980 32525
rect 14600 32925 14736 32966
rect 14600 32567 14680 32925
rect 14723 32787 14781 32790
rect 14723 32735 14726 32787
rect 14778 32735 14781 32787
rect 14723 32732 14781 32735
rect 14600 32525 14736 32567
rect 14600 32218 14680 32525
rect 14723 32387 14781 32390
rect 14723 32335 14726 32387
rect 14778 32335 14781 32387
rect 14723 32332 14781 32335
rect 4900 32167 4951 32218
rect 4844 32166 4951 32167
rect 4977 32166 4980 32218
rect 14600 32166 14603 32218
rect 14629 32167 14680 32218
rect 14629 32166 14736 32167
rect 4844 32125 4980 32166
rect 4799 31987 4857 31990
rect 4799 31935 4802 31987
rect 4854 31935 4857 31987
rect 4799 31932 4857 31935
rect 4900 31767 4980 32125
rect 4844 31725 4980 31767
rect 4799 31587 4857 31590
rect 4799 31535 4802 31587
rect 4854 31535 4857 31587
rect 4799 31532 4857 31535
rect 4900 31418 4980 31725
rect 14600 32125 14736 32166
rect 14600 31767 14680 32125
rect 14723 31987 14781 31990
rect 14723 31935 14726 31987
rect 14778 31935 14781 31987
rect 14723 31932 14781 31935
rect 14600 31725 14736 31767
rect 14600 31418 14680 31725
rect 14723 31587 14781 31590
rect 14723 31535 14726 31587
rect 14778 31535 14781 31587
rect 14723 31532 14781 31535
rect 4900 31367 4951 31418
rect 4844 31366 4951 31367
rect 4977 31366 4980 31418
rect 14600 31366 14603 31418
rect 14629 31367 14680 31418
rect 14629 31366 14736 31367
rect 4844 31325 4980 31366
rect 4799 31187 4857 31190
rect 4799 31135 4802 31187
rect 4854 31135 4857 31187
rect 4799 31132 4857 31135
rect 4900 30967 4980 31325
rect 4844 30925 4980 30967
rect 4799 30787 4857 30790
rect 4799 30735 4802 30787
rect 4854 30735 4857 30787
rect 4799 30732 4857 30735
rect 4900 30618 4980 30925
rect 14600 31325 14736 31366
rect 14600 30967 14680 31325
rect 14723 31187 14781 31190
rect 14723 31135 14726 31187
rect 14778 31135 14781 31187
rect 14723 31132 14781 31135
rect 14600 30925 14736 30967
rect 14600 30618 14680 30925
rect 14723 30787 14781 30790
rect 14723 30735 14726 30787
rect 14778 30735 14781 30787
rect 14723 30732 14781 30735
rect 4900 30567 4951 30618
rect 4844 30566 4951 30567
rect 4977 30566 4980 30618
rect 14600 30566 14603 30618
rect 14629 30567 14680 30618
rect 14629 30566 14736 30567
rect 4844 30525 4980 30566
rect 4799 30387 4857 30390
rect 4799 30335 4802 30387
rect 4854 30335 4857 30387
rect 4799 30332 4857 30335
rect 4900 30167 4980 30525
rect 4844 30125 4980 30167
rect 4799 29987 4857 29990
rect 4799 29935 4802 29987
rect 4854 29935 4857 29987
rect 4799 29932 4857 29935
rect 4900 29818 4980 30125
rect 14600 30525 14736 30566
rect 14600 30167 14680 30525
rect 14723 30387 14781 30390
rect 14723 30335 14726 30387
rect 14778 30335 14781 30387
rect 14723 30332 14781 30335
rect 14600 30125 14736 30167
rect 14600 29818 14680 30125
rect 14723 29987 14781 29990
rect 14723 29935 14726 29987
rect 14778 29935 14781 29987
rect 14723 29932 14781 29935
rect 4900 29767 4951 29818
rect 4844 29766 4951 29767
rect 4977 29766 4980 29818
rect 14600 29766 14603 29818
rect 14629 29767 14680 29818
rect 14629 29766 14736 29767
rect 4844 29725 4980 29766
rect 4799 29587 4857 29590
rect 4799 29535 4802 29587
rect 4854 29535 4857 29587
rect 4799 29532 4857 29535
rect 4900 29367 4980 29725
rect 4844 29325 4980 29367
rect 14600 29725 14736 29766
rect 14600 29367 14680 29725
rect 14723 29587 14781 29590
rect 14723 29535 14726 29587
rect 14778 29535 14781 29587
rect 14723 29532 14781 29535
rect 14600 29325 14736 29367
rect 4799 29187 4857 29190
rect 4799 29135 4802 29187
rect 4854 29135 4857 29187
rect 4799 29132 4857 29135
rect 14723 29187 14781 29190
rect 14723 29135 14726 29187
rect 14778 29135 14781 29187
rect 14723 29132 14781 29135
<< via1 >>
rect 4900 41793 4980 41871
rect 14600 41793 14680 41871
rect 4802 41535 4854 41587
rect 4802 41135 4854 41187
rect 14726 41535 14778 41587
rect 14726 41135 14778 41187
rect 4951 40966 4977 41018
rect 5130 40966 5156 41018
rect 14424 40966 14450 41018
rect 14603 40966 14629 41018
rect 4802 40735 4854 40787
rect 4802 40335 4854 40387
rect 14726 40735 14778 40787
rect 14726 40335 14778 40387
rect 4951 40166 4977 40218
rect 5130 40166 5156 40218
rect 14424 40166 14450 40218
rect 14603 40166 14629 40218
rect 4802 39935 4854 39987
rect 4802 39535 4854 39587
rect 14726 39935 14778 39987
rect 14726 39535 14778 39587
rect 4951 39366 4977 39418
rect 5130 39366 5156 39418
rect 14424 39366 14450 39418
rect 14603 39366 14629 39418
rect 4802 39135 4854 39187
rect 4802 38735 4854 38787
rect 14726 39135 14778 39187
rect 14726 38735 14778 38787
rect 4951 38566 4977 38618
rect 5130 38566 5156 38618
rect 14424 38566 14450 38618
rect 14603 38566 14629 38618
rect 4802 38335 4854 38387
rect 4802 37935 4854 37987
rect 14726 38335 14778 38387
rect 14726 37935 14778 37987
rect 4951 37766 4977 37818
rect 5130 37766 5156 37818
rect 14424 37766 14450 37818
rect 14603 37766 14629 37818
rect 4802 37535 4854 37587
rect 4802 37135 4854 37187
rect 14726 37535 14778 37587
rect 14726 37135 14778 37187
rect 4951 36966 4977 37018
rect 5130 36966 5156 37018
rect 14424 36966 14450 37018
rect 14603 36966 14629 37018
rect 4802 36735 4854 36787
rect 4802 36335 4854 36387
rect 14726 36735 14778 36787
rect 14726 36335 14778 36387
rect 4951 36166 4977 36218
rect 5130 36166 5156 36218
rect 14424 36166 14450 36218
rect 14603 36166 14629 36218
rect 4802 35935 4854 35987
rect 4802 35535 4854 35587
rect 14726 35935 14778 35987
rect 14726 35535 14778 35587
rect 4951 35366 4977 35418
rect 5130 35366 5156 35418
rect 14424 35366 14450 35418
rect 14603 35366 14629 35418
rect 4802 35135 4854 35187
rect 4802 34735 4854 34787
rect 14726 35135 14778 35187
rect 14726 34735 14778 34787
rect 4951 34566 4977 34618
rect 5130 34566 5156 34618
rect 14424 34566 14450 34618
rect 14603 34566 14629 34618
rect 4802 34335 4854 34387
rect 4802 33935 4854 33987
rect 14726 34335 14778 34387
rect 14726 33935 14778 33987
rect 4951 33766 4977 33818
rect 5130 33766 5156 33818
rect 14424 33766 14450 33818
rect 14603 33766 14629 33818
rect 4802 33535 4854 33587
rect 4802 33135 4854 33187
rect 14726 33535 14778 33587
rect 14726 33135 14778 33187
rect 4951 32966 4977 33018
rect 5130 32966 5156 33018
rect 14424 32966 14450 33018
rect 14603 32966 14629 33018
rect 4802 32735 4854 32787
rect 4802 32335 4854 32387
rect 14726 32735 14778 32787
rect 14726 32335 14778 32387
rect 4951 32166 4977 32218
rect 5130 32166 5156 32218
rect 14424 32166 14450 32218
rect 14603 32166 14629 32218
rect 4802 31935 4854 31987
rect 4802 31535 4854 31587
rect 14726 31935 14778 31987
rect 14726 31535 14778 31587
rect 4951 31366 4977 31418
rect 5130 31366 5156 31418
rect 14424 31366 14450 31418
rect 14603 31366 14629 31418
rect 4802 31135 4854 31187
rect 4802 30735 4854 30787
rect 14726 31135 14778 31187
rect 14726 30735 14778 30787
rect 4951 30566 4977 30618
rect 5130 30566 5156 30618
rect 14424 30566 14450 30618
rect 14603 30566 14629 30618
rect 4802 30335 4854 30387
rect 4802 29935 4854 29987
rect 14726 30335 14778 30387
rect 14726 29935 14778 29987
rect 4951 29766 4977 29818
rect 5130 29766 5156 29818
rect 14424 29766 14450 29818
rect 14603 29766 14629 29818
rect 4802 29535 4854 29587
rect 14726 29535 14778 29587
rect 4802 29135 4854 29187
rect 14726 29135 14778 29187
<< metal2 >>
rect 4897 41793 4900 41871
rect 4980 41793 5130 41871
rect 14450 41793 14600 41871
rect 14680 41793 14683 41871
rect 4799 41587 5000 41590
rect 4799 41535 4802 41587
rect 4854 41535 5000 41587
rect 4799 41532 5000 41535
rect 14580 41587 14781 41590
rect 14580 41535 14726 41587
rect 14778 41535 14781 41587
rect 14580 41532 14781 41535
rect 4799 41187 5000 41190
rect 4799 41135 4802 41187
rect 4854 41135 5000 41187
rect 4799 41132 5000 41135
rect 14580 41187 14781 41190
rect 14580 41135 14726 41187
rect 14778 41135 14781 41187
rect 14580 41132 14781 41135
rect 4948 41018 5159 41021
rect 4948 40966 4951 41018
rect 4977 40966 5130 41018
rect 5156 40966 5159 41018
rect 4948 40963 5159 40966
rect 14421 41018 14632 41021
rect 14421 40966 14424 41018
rect 14450 40966 14603 41018
rect 14629 40966 14632 41018
rect 14421 40963 14632 40966
rect 4799 40787 5000 40790
rect 4799 40735 4802 40787
rect 4854 40735 5000 40787
rect 4799 40732 5000 40735
rect 14580 40787 14781 40790
rect 14580 40735 14726 40787
rect 14778 40735 14781 40787
rect 14580 40732 14781 40735
rect 4799 40387 5000 40390
rect 4799 40335 4802 40387
rect 4854 40335 5000 40387
rect 4799 40332 5000 40335
rect 14580 40387 14781 40390
rect 14580 40335 14726 40387
rect 14778 40335 14781 40387
rect 14580 40332 14781 40335
rect 4948 40218 5159 40221
rect 4948 40166 4951 40218
rect 4977 40166 5130 40218
rect 5156 40166 5159 40218
rect 4948 40163 5159 40166
rect 14421 40218 14632 40221
rect 14421 40166 14424 40218
rect 14450 40166 14603 40218
rect 14629 40166 14632 40218
rect 14421 40163 14632 40166
rect 4799 39987 5000 39990
rect 4799 39935 4802 39987
rect 4854 39935 5000 39987
rect 4799 39932 5000 39935
rect 14580 39987 14781 39990
rect 14580 39935 14726 39987
rect 14778 39935 14781 39987
rect 14580 39932 14781 39935
rect 4799 39587 5000 39590
rect 4799 39535 4802 39587
rect 4854 39535 5000 39587
rect 4799 39532 5000 39535
rect 14580 39587 14781 39590
rect 14580 39535 14726 39587
rect 14778 39535 14781 39587
rect 14580 39532 14781 39535
rect 4948 39418 5159 39421
rect 4948 39366 4951 39418
rect 4977 39366 5130 39418
rect 5156 39366 5159 39418
rect 4948 39363 5159 39366
rect 14421 39418 14632 39421
rect 14421 39366 14424 39418
rect 14450 39366 14603 39418
rect 14629 39366 14632 39418
rect 14421 39363 14632 39366
rect 4799 39187 5000 39190
rect 4799 39135 4802 39187
rect 4854 39135 5000 39187
rect 4799 39132 5000 39135
rect 14580 39187 14781 39190
rect 14580 39135 14726 39187
rect 14778 39135 14781 39187
rect 14580 39132 14781 39135
rect 4799 38787 5000 38790
rect 4799 38735 4802 38787
rect 4854 38735 5000 38787
rect 4799 38732 5000 38735
rect 14580 38787 14781 38790
rect 14580 38735 14726 38787
rect 14778 38735 14781 38787
rect 14580 38732 14781 38735
rect 4948 38618 5159 38621
rect 4948 38566 4951 38618
rect 4977 38566 5130 38618
rect 5156 38566 5159 38618
rect 4948 38563 5159 38566
rect 14421 38618 14632 38621
rect 14421 38566 14424 38618
rect 14450 38566 14603 38618
rect 14629 38566 14632 38618
rect 14421 38563 14632 38566
rect 4799 38387 5000 38390
rect 4799 38335 4802 38387
rect 4854 38335 5000 38387
rect 4799 38332 5000 38335
rect 14580 38387 14781 38390
rect 14580 38335 14726 38387
rect 14778 38335 14781 38387
rect 14580 38332 14781 38335
rect 4799 37987 5000 37990
rect 4799 37935 4802 37987
rect 4854 37935 5000 37987
rect 4799 37932 5000 37935
rect 14580 37987 14781 37990
rect 14580 37935 14726 37987
rect 14778 37935 14781 37987
rect 14580 37932 14781 37935
rect 4948 37818 5159 37821
rect 4948 37766 4951 37818
rect 4977 37766 5130 37818
rect 5156 37766 5159 37818
rect 4948 37763 5159 37766
rect 14421 37818 14632 37821
rect 14421 37766 14424 37818
rect 14450 37766 14603 37818
rect 14629 37766 14632 37818
rect 14421 37763 14632 37766
rect 4799 37587 5000 37590
rect 4799 37535 4802 37587
rect 4854 37535 5000 37587
rect 4799 37532 5000 37535
rect 14580 37587 14781 37590
rect 14580 37535 14726 37587
rect 14778 37535 14781 37587
rect 14580 37532 14781 37535
rect 4799 37187 5000 37190
rect 4799 37135 4802 37187
rect 4854 37135 5000 37187
rect 4799 37132 5000 37135
rect 14580 37187 14781 37190
rect 14580 37135 14726 37187
rect 14778 37135 14781 37187
rect 14580 37132 14781 37135
rect 4948 37018 5159 37021
rect 4948 36966 4951 37018
rect 4977 36966 5130 37018
rect 5156 36966 5159 37018
rect 4948 36963 5159 36966
rect 14421 37018 14632 37021
rect 14421 36966 14424 37018
rect 14450 36966 14603 37018
rect 14629 36966 14632 37018
rect 14421 36963 14632 36966
rect 4799 36787 5000 36790
rect 4799 36735 4802 36787
rect 4854 36735 5000 36787
rect 4799 36732 5000 36735
rect 14580 36787 14781 36790
rect 14580 36735 14726 36787
rect 14778 36735 14781 36787
rect 14580 36732 14781 36735
rect 4799 36387 5000 36390
rect 4799 36335 4802 36387
rect 4854 36335 5000 36387
rect 4799 36332 5000 36335
rect 14580 36387 14781 36390
rect 14580 36335 14726 36387
rect 14778 36335 14781 36387
rect 14580 36332 14781 36335
rect 4948 36218 5159 36221
rect 4948 36166 4951 36218
rect 4977 36166 5130 36218
rect 5156 36166 5159 36218
rect 4948 36163 5159 36166
rect 14421 36218 14632 36221
rect 14421 36166 14424 36218
rect 14450 36166 14603 36218
rect 14629 36166 14632 36218
rect 14421 36163 14632 36166
rect 4799 35987 5000 35990
rect 4799 35935 4802 35987
rect 4854 35935 5000 35987
rect 4799 35932 5000 35935
rect 14580 35987 14781 35990
rect 14580 35935 14726 35987
rect 14778 35935 14781 35987
rect 14580 35932 14781 35935
rect 4799 35587 5000 35590
rect 4799 35535 4802 35587
rect 4854 35535 5000 35587
rect 4799 35532 5000 35535
rect 14580 35587 14781 35590
rect 14580 35535 14726 35587
rect 14778 35535 14781 35587
rect 14580 35532 14781 35535
rect 4948 35418 5159 35421
rect 4948 35366 4951 35418
rect 4977 35366 5130 35418
rect 5156 35366 5159 35418
rect 4948 35363 5159 35366
rect 14421 35418 14632 35421
rect 14421 35366 14424 35418
rect 14450 35366 14603 35418
rect 14629 35366 14632 35418
rect 14421 35363 14632 35366
rect 4799 35187 5000 35190
rect 4799 35135 4802 35187
rect 4854 35135 5000 35187
rect 4799 35132 5000 35135
rect 14580 35187 14781 35190
rect 14580 35135 14726 35187
rect 14778 35135 14781 35187
rect 14580 35132 14781 35135
rect 4799 34787 5000 34790
rect 4799 34735 4802 34787
rect 4854 34735 5000 34787
rect 4799 34732 5000 34735
rect 14580 34787 14781 34790
rect 14580 34735 14726 34787
rect 14778 34735 14781 34787
rect 14580 34732 14781 34735
rect 4948 34618 5159 34621
rect 4948 34566 4951 34618
rect 4977 34566 5130 34618
rect 5156 34566 5159 34618
rect 4948 34563 5159 34566
rect 14421 34618 14632 34621
rect 14421 34566 14424 34618
rect 14450 34566 14603 34618
rect 14629 34566 14632 34618
rect 14421 34563 14632 34566
rect 4799 34387 5000 34390
rect 4799 34335 4802 34387
rect 4854 34335 5000 34387
rect 4799 34332 5000 34335
rect 14580 34387 14781 34390
rect 14580 34335 14726 34387
rect 14778 34335 14781 34387
rect 14580 34332 14781 34335
rect 4799 33987 5000 33990
rect 4799 33935 4802 33987
rect 4854 33935 5000 33987
rect 4799 33932 5000 33935
rect 14580 33987 14781 33990
rect 14580 33935 14726 33987
rect 14778 33935 14781 33987
rect 14580 33932 14781 33935
rect 4948 33818 5159 33821
rect 4948 33766 4951 33818
rect 4977 33766 5130 33818
rect 5156 33766 5159 33818
rect 4948 33763 5159 33766
rect 14421 33818 14632 33821
rect 14421 33766 14424 33818
rect 14450 33766 14603 33818
rect 14629 33766 14632 33818
rect 14421 33763 14632 33766
rect 4799 33587 5000 33590
rect 4799 33535 4802 33587
rect 4854 33535 5000 33587
rect 4799 33532 5000 33535
rect 14580 33587 14781 33590
rect 14580 33535 14726 33587
rect 14778 33535 14781 33587
rect 14580 33532 14781 33535
rect 4799 33187 5000 33190
rect 4799 33135 4802 33187
rect 4854 33135 5000 33187
rect 4799 33132 5000 33135
rect 14580 33187 14781 33190
rect 14580 33135 14726 33187
rect 14778 33135 14781 33187
rect 14580 33132 14781 33135
rect 4948 33018 5159 33021
rect 4948 32966 4951 33018
rect 4977 32966 5130 33018
rect 5156 32966 5159 33018
rect 4948 32963 5159 32966
rect 14421 33018 14632 33021
rect 14421 32966 14424 33018
rect 14450 32966 14603 33018
rect 14629 32966 14632 33018
rect 14421 32963 14632 32966
rect 4799 32787 5000 32790
rect 4799 32735 4802 32787
rect 4854 32735 5000 32787
rect 4799 32732 5000 32735
rect 14580 32787 14781 32790
rect 14580 32735 14726 32787
rect 14778 32735 14781 32787
rect 14580 32732 14781 32735
rect 4799 32387 5000 32390
rect 4799 32335 4802 32387
rect 4854 32335 5000 32387
rect 4799 32332 5000 32335
rect 14580 32387 14781 32390
rect 14580 32335 14726 32387
rect 14778 32335 14781 32387
rect 14580 32332 14781 32335
rect 4948 32218 5159 32221
rect 4948 32166 4951 32218
rect 4977 32166 5130 32218
rect 5156 32166 5159 32218
rect 4948 32163 5159 32166
rect 14421 32218 14632 32221
rect 14421 32166 14424 32218
rect 14450 32166 14603 32218
rect 14629 32166 14632 32218
rect 14421 32163 14632 32166
rect 4799 31987 5000 31990
rect 4799 31935 4802 31987
rect 4854 31935 5000 31987
rect 4799 31932 5000 31935
rect 14580 31987 14781 31990
rect 14580 31935 14726 31987
rect 14778 31935 14781 31987
rect 14580 31932 14781 31935
rect 4799 31587 5000 31590
rect 4799 31535 4802 31587
rect 4854 31535 5000 31587
rect 4799 31532 5000 31535
rect 14580 31587 14781 31590
rect 14580 31535 14726 31587
rect 14778 31535 14781 31587
rect 14580 31532 14781 31535
rect 4948 31418 5159 31421
rect 4948 31366 4951 31418
rect 4977 31366 5130 31418
rect 5156 31366 5159 31418
rect 4948 31363 5159 31366
rect 14421 31418 14632 31421
rect 14421 31366 14424 31418
rect 14450 31366 14603 31418
rect 14629 31366 14632 31418
rect 14421 31363 14632 31366
rect 4799 31187 5000 31190
rect 4799 31135 4802 31187
rect 4854 31135 5000 31187
rect 4799 31132 5000 31135
rect 14580 31187 14781 31190
rect 14580 31135 14726 31187
rect 14778 31135 14781 31187
rect 14580 31132 14781 31135
rect 4799 30787 5000 30790
rect 4799 30735 4802 30787
rect 4854 30735 5000 30787
rect 4799 30732 5000 30735
rect 14580 30787 14781 30790
rect 14580 30735 14726 30787
rect 14778 30735 14781 30787
rect 14580 30732 14781 30735
rect 4948 30618 5159 30621
rect 4948 30566 4951 30618
rect 4977 30566 5130 30618
rect 5156 30566 5159 30618
rect 4948 30563 5159 30566
rect 14421 30618 14632 30621
rect 14421 30566 14424 30618
rect 14450 30566 14603 30618
rect 14629 30566 14632 30618
rect 14421 30563 14632 30566
rect 4799 30387 5000 30390
rect 4799 30335 4802 30387
rect 4854 30335 5000 30387
rect 4799 30332 5000 30335
rect 14580 30387 14781 30390
rect 14580 30335 14726 30387
rect 14778 30335 14781 30387
rect 14580 30332 14781 30335
rect 4799 29987 5000 29990
rect 4799 29935 4802 29987
rect 4854 29935 5000 29987
rect 4799 29932 5000 29935
rect 14580 29987 14781 29990
rect 14580 29935 14726 29987
rect 14778 29935 14781 29987
rect 14580 29932 14781 29935
rect 4948 29818 5159 29821
rect 4948 29766 4951 29818
rect 4977 29766 5130 29818
rect 5156 29766 5159 29818
rect 4948 29763 5159 29766
rect 14421 29818 14632 29821
rect 14421 29766 14424 29818
rect 14450 29766 14603 29818
rect 14629 29766 14632 29818
rect 14421 29763 14632 29766
rect 4799 29587 5000 29590
rect 4799 29535 4802 29587
rect 4854 29535 5000 29587
rect 4799 29532 5000 29535
rect 14580 29587 14781 29590
rect 14580 29535 14726 29587
rect 14778 29535 14781 29587
rect 14580 29532 14781 29535
rect 4799 29187 5000 29190
rect 4799 29135 4802 29187
rect 4854 29135 5000 29187
rect 4799 29132 5000 29135
rect 14580 29187 14781 29190
rect 14580 29135 14726 29187
rect 14778 29135 14781 29187
rect 14580 29132 14781 29135
use array_core_block0  array_core_block0_0
timestamp 1717164735
transform 1 0 -20000 0 1 30696
box 0 -696 19983 14118
use array_core_block1  array_core_block1_0
timestamp 1717164735
transform 1 0 -20000 0 1 15000
box 0 0 19983 14814
use array_core_block2  array_core_block2_0
timestamp 1717164735
transform 1 0 -20000 0 1 0
box 0 0 19983 14819
use array_core_block3  array_core_block3_0
timestamp 1717164735
transform 1 0 20000 0 1 30000
box 0 0 19983 14411
use array_core_block4  array_core_block4_0
timestamp 1717164735
transform 1 0 20000 0 1 15000
box 0 0 19983 14411
use array_core_block5  array_core_block5_0
timestamp 1717164252
transform 1 0 20033 0 1 0
box -33 0 19983 14623
use array_row_decode  array_row_decode_0
timestamp 1717093521
transform 1 0 13020 0 1 28832
box -2020 168 1560 14074
use array_row_decode  array_row_decode_1
timestamp 1717093521
transform -1 0 6560 0 1 28832
box -2020 168 1560 14074
use lsi1v8o5v0  lsi1v8o5v0_0
array 0 0 1161 0 31 -400
timestamp 1717165718
transform -1 0 4858 0 -1 29307
box -42 -60 1119 293
use lsi1v8o5v0  lsi1v8o5v0_1
array 0 0 1161 0 31 -400
timestamp 1717165718
transform 1 0 14722 0 -1 29307
box -42 -60 1119 293
<< end >>
