magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< error_s >>
rect 2122 -5050 2442 -4988
rect 506 -5294 746 -5270
rect 506 -5486 530 -5294
rect 722 -5486 746 -5294
rect 2122 -5290 2146 -5050
rect 2382 -5290 2386 -5050
rect 2406 -5290 2442 -5050
rect 2122 -5314 2442 -5290
rect 506 -5510 746 -5486
rect 2996 -5499 3132 -5494
rect 2996 -5573 3001 -5499
rect 3127 -5573 3132 -5499
rect 2996 -5578 3132 -5573
rect 2506 -5651 2686 -5650
rect 2506 -5829 2507 -5651
rect 2685 -5829 2686 -5651
rect 2506 -5830 2686 -5829
rect 3868 -6200 3874 -6194
rect 3920 -6200 3926 -6194
rect 3862 -6206 3868 -6200
rect 3926 -6206 3932 -6200
rect 526 -6211 706 -6210
rect 526 -6389 527 -6211
rect 705 -6389 706 -6211
rect 3862 -6262 3868 -6256
rect 3926 -6262 3932 -6256
rect 3868 -6268 3874 -6262
rect 3920 -6268 3926 -6262
rect 526 -6390 706 -6389
rect 3402 -6402 3408 -6396
rect 3448 -6402 3454 -6396
rect 3396 -6408 3402 -6402
rect 3454 -6408 3460 -6402
rect 3396 -6454 3402 -6448
rect 3454 -6454 3460 -6448
rect 3402 -6460 3408 -6454
rect 3448 -6460 3454 -6454
rect 2426 -6914 2666 -6890
rect 2426 -7106 2450 -6914
rect 2642 -7106 2666 -6914
rect 2426 -7130 2666 -7106
<< mvnmos >>
rect 1336 -5964 2938 -5864
<< mvndiff >>
rect 1282 -5864 2938 -5814
rect 1282 -5964 1336 -5864
rect 1282 -6014 2938 -5964
<< poly >>
rect 2907 -5477 3240 -5380
rect 3140 -5864 3240 -5477
rect 2938 -5964 3240 -5864
rect 3140 -6470 3240 -5964
<< locali >>
rect 3076 -5190 3282 -5060
<< metal1 >>
rect 2126 -5050 2406 -5030
rect 2126 -5290 2146 -5050
rect 2386 -5290 2406 -5050
rect 2496 -5050 2656 -5040
rect 2496 -5190 2506 -5050
rect 2646 -5190 2656 -5050
rect 3736 -5042 3836 -5036
rect 3076 -5190 3322 -5098
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3736 -5130 3742 -5042
rect 3830 -5130 3836 -5042
rect 3736 -5136 3836 -5130
rect 2496 -5198 2656 -5190
rect 3360 -5194 3460 -5188
rect 2126 -5310 2406 -5290
rect 3868 -6200 3932 -6194
rect 3926 -6262 3932 -6200
rect 3868 -6268 3932 -6262
rect 3868 -6384 3872 -6378
rect 3396 -6402 3454 -6396
rect 3396 -6454 3402 -6402
rect 3396 -6458 3454 -6454
rect 3868 -6458 3872 -6446
rect 3134 -6806 3240 -6570
rect 3502 -6806 3604 -6558
rect 3134 -6812 3604 -6806
rect 3134 -6900 3140 -6812
rect 3234 -6900 3604 -6812
rect 3134 -6904 3604 -6900
rect 3134 -6906 3240 -6904
rect 2476 -7030 2676 -7020
rect 4006 -7030 4106 -5098
rect 2476 -7130 2486 -7030
rect 2666 -7130 2676 -7030
rect 2900 -7130 4106 -7030
rect 2476 -7140 2676 -7130
<< via1 >>
rect 2146 -5290 2386 -5050
rect 2506 -5190 2646 -5050
rect 3366 -5188 3454 -5100
rect 3742 -5130 3830 -5042
rect 3868 -6262 3926 -6200
rect 3402 -6454 3454 -6402
rect 3140 -6900 3234 -6812
rect 406 -7104 914 -7036
rect 2486 -7130 2666 -7030
<< metal2 >>
rect 2126 -5050 2406 -5030
rect 506 -5270 746 -5260
rect 2126 -5290 2146 -5050
rect 2386 -5290 2406 -5050
rect 2496 -5050 2656 -5040
rect 2496 -5190 2506 -5050
rect 2646 -5190 2656 -5050
rect 3732 -5042 3840 -5032
rect 2496 -5200 2656 -5190
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3732 -5130 3742 -5042
rect 3830 -5130 3840 -5042
rect 3732 -5140 3840 -5130
rect 3360 -5222 3460 -5188
rect 2126 -5310 2406 -5290
rect 2938 -5322 3460 -5222
rect 506 -5520 746 -5510
rect 2758 -5494 3142 -5484
rect 2758 -5578 2996 -5494
rect 3132 -5578 3142 -5494
rect 2758 -5588 3142 -5578
rect 1294 -6812 3240 -6806
rect 1294 -6900 3140 -6812
rect 3234 -6900 3240 -6812
rect 1294 -6906 3240 -6900
rect 520 -6924 712 -6914
rect 520 -7030 526 -6924
rect 396 -7036 526 -7030
rect 706 -7030 712 -6924
rect 2476 -7030 2676 -7020
rect 706 -7036 924 -7030
rect 396 -7104 406 -7036
rect 914 -7104 924 -7036
rect 396 -7110 924 -7104
rect 520 -7114 712 -7110
rect 2476 -7130 2486 -7030
rect 2666 -7130 2676 -7030
rect 2476 -7140 2676 -7130
<< via2 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2506 -5190 2646 -5050
rect 3742 -5130 3830 -5042
rect 2996 -5578 3132 -5494
rect 526 -7036 706 -6924
rect 526 -7104 706 -7036
rect 2486 -7130 2666 -7030
<< metal3 >>
rect 2126 -5050 2406 -5030
rect 500 -5270 752 -5264
rect 500 -5510 506 -5270
rect 746 -5510 752 -5270
rect 2126 -5290 2146 -5050
rect 2386 -5290 2406 -5050
rect 2126 -5310 2406 -5290
rect 2486 -5050 2706 -5030
rect 2486 -5190 2506 -5050
rect 2646 -5190 2706 -5050
rect 3732 -5042 3840 -5032
rect 3732 -5130 3742 -5042
rect 3830 -5130 3840 -5042
rect 3732 -5140 3840 -5130
rect 500 -5516 752 -5510
rect 2486 -5650 2706 -5190
rect 2486 -5830 2506 -5650
rect 2686 -5830 2706 -5650
rect 2486 -5850 2706 -5830
rect 520 -6210 712 -6204
rect 520 -6390 526 -6210
rect 706 -6390 712 -6210
rect 520 -6924 712 -6390
rect 520 -7104 526 -6924
rect 706 -7104 712 -6924
rect 520 -7110 712 -7104
rect 2422 -6950 2676 -6886
rect 2422 -7130 2486 -6950
rect 2666 -7130 2676 -6950
rect 2422 -7140 2676 -7130
<< via3 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2506 -5830 2686 -5650
rect 526 -6390 706 -6210
rect 2486 -7030 2666 -6950
rect 2486 -7130 2666 -7030
<< metal4 >>
rect 2126 -5050 2406 -5030
rect 500 -5270 752 -5264
rect 500 -5510 506 -5270
rect 746 -5510 752 -5270
rect 2126 -5290 2146 -5050
rect 2386 -5290 2406 -5050
rect 2126 -5314 2406 -5290
rect 500 -5516 752 -5510
rect 2422 -6890 2676 -6886
rect 2422 -7130 2426 -6890
rect 2666 -7130 2676 -6890
rect 2422 -7140 2676 -7130
<< via4 >>
rect 506 -5510 746 -5270
rect 2146 -5290 2386 -5050
rect 2426 -6950 2666 -6890
rect 2426 -7130 2486 -6950
rect 2486 -7130 2666 -6950
<< metal5 >>
rect 2122 -5050 2406 -4988
rect 2122 -5290 2146 -5050
rect 2386 -5290 2406 -5050
rect 2122 -5314 2406 -5290
use tg5v0  tg5v0_0
timestamp 1717628967
transform 0 -1 4094 1 0 -6628
box 28 0 1634 890
use fgcell  x1
timestamp 1717628967
transform 1 0 2010 0 1 -5490
box -1870 -310 1194 526
use diffamp_nmos  x2
timestamp 1717628967
transform 0 -1 3100 -1 0 -6070
box 20 -140 1140 2900
<< labels >>
flabel via2 2996 -5578 3132 -5494 0 FreeSans 320 0 0 0 vsrc
flabel via4 2146 -5290 2386 -5050 0 FreeSans 320 0 0 0 VGND
flabel via4 2426 -7130 2666 -6890 0 FreeSans 320 0 0 0 VGND
flabel via4 506 -5510 746 -5270 0 FreeSans 320 0 0 0 vtun
flabel via3 526 -6390 706 -6210 0 FreeSans 640 0 0 0 vdd
flabel via1 3402 -6454 3454 -6402 0 FreeSans 32 0 0 0 row_en_b
flabel via1 3868 -6262 3926 -6200 0 FreeSans 320 0 0 0 row_en
<< end >>
