** sch_path: /home/amedcalf/projects/ci2406_fgcaptest/xschem/tb_diffamp_nmos_ac.sch
**.subckt tb_diffamp_nmos_ac
x1 v1 vout GND VDD vb vout diffamp_nmos
VDD VDD GND {VDD}
vb vb GND {VBIAS}
v1 v1 GND dc 3 ac 1 sin(3 1 1meg)
R1 vout GND 1g m=1
v2 net1 GND 3
C1 vout GND 26f m=1
**** begin user architecture code
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.options reltol=0.0001 abstol=10e-15
.include diffamp_nmos.spice
.param VDD=5
.param VSS=0
.param VBIAS=1
.options savecurrents
* .options reltol=0.01 abstol=10e-12
.control
  save all
  op
  remzerovec
  write tb_diffamp_nmos_ac.raw
  set appendwrite
  * ac sweep
  ac dec 20 1 1gig
  remzerovec
  write tb_diffamp_nmos_ac.raw
  * tran
  tran 1n 5u
  remzerovec
  write tb_diffamp_nmos_ac.raw
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
