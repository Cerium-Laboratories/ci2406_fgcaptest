magic
tech sky130A
magscale 1 2
timestamp 1716414739
<< nwell >>
rect -1576 -75 -1194 291
rect -710 -200 -84 416
rect 400 -248 1194 526
<< mvpmos >>
rect 697 168 897 268
rect -497 58 -297 158
rect 697 10 897 110
<< varactorhvt >>
rect -1485 58 -1285 158
<< mvpdiff >>
rect 697 314 897 326
rect 697 280 709 314
rect 885 280 897 314
rect 697 268 897 280
rect -497 204 -297 216
rect -497 170 -485 204
rect -309 170 -297 204
rect -497 158 -297 170
rect 697 110 897 168
rect -497 46 -297 58
rect -497 12 -485 46
rect -309 12 -297 46
rect -497 0 -297 12
rect 697 -2 897 10
rect 697 -36 709 -2
rect 885 -36 897 -2
rect 697 -48 897 -36
<< mvpdiffc >>
rect 709 280 885 314
rect -485 170 -309 204
rect -485 12 -309 46
rect 709 -36 885 -2
<< psubdiff >>
rect -1810 506 -960 526
rect -1810 466 -1730 506
rect -1040 466 -960 506
rect -1810 446 -960 466
rect -1810 392 -1730 446
rect -1810 -176 -1790 392
rect -1750 -176 -1730 392
rect -1040 392 -960 446
rect -1040 252 -1020 392
rect -980 252 -960 392
rect 160 392 240 416
rect -1040 228 -960 252
rect 160 252 180 392
rect 220 252 240 392
rect 160 228 240 252
rect -1040 -36 -960 -12
rect -1810 -230 -1730 -176
rect -1040 -176 -1020 -36
rect -980 -176 -960 -36
rect 160 -36 240 -12
rect -1040 -230 -960 -176
rect 160 -176 180 -36
rect 220 -176 240 -36
rect 160 -200 240 -176
rect -1810 -250 -960 -230
rect -1810 -290 -1730 -250
rect -1040 -290 -960 -250
rect -1810 -310 -960 -290
<< nsubdiff >>
rect -1485 243 -1285 255
rect -1485 209 -1461 243
rect -1309 209 -1285 243
rect -1485 158 -1285 209
rect -1485 7 -1285 58
rect -1485 -27 -1461 7
rect -1309 -27 -1285 7
rect -1485 -39 -1285 -27
<< mvnsubdiff >>
rect 466 448 1128 460
rect 466 414 574 448
rect 1020 414 1128 448
rect 466 402 1128 414
rect -644 338 -150 350
rect -644 304 -620 338
rect -174 304 -150 338
rect -644 292 -150 304
rect 1070 352 1128 402
rect 1070 194 1082 352
rect 1116 194 1128 352
rect 1070 84 1128 194
rect -644 -88 -150 -76
rect -644 -122 -620 -88
rect -174 -122 -150 -88
rect -644 -134 -150 -122
rect 1070 -74 1082 84
rect 1116 -74 1128 84
rect 1070 -124 1128 -74
rect 466 -136 1128 -124
rect 466 -170 574 -136
rect 1020 -170 1128 -136
rect 466 -182 1128 -170
<< psubdiffcont >>
rect -1730 466 -1040 506
rect -1790 -176 -1750 392
rect -1020 252 -980 392
rect 180 252 220 392
rect -1020 -176 -980 -36
rect 180 -176 220 -36
rect -1730 -290 -1040 -250
<< nsubdiffcont >>
rect -1461 209 -1309 243
rect -1461 -27 -1309 7
<< mvnsubdiffcont >>
rect 574 414 1020 448
rect -620 304 -174 338
rect 1082 194 1116 352
rect -620 -122 -174 -88
rect 1082 -74 1116 84
rect 574 -170 1020 -136
<< poly >>
rect 600 252 697 268
rect 600 184 616 252
rect 650 184 697 252
rect 600 168 697 184
rect 897 168 994 268
rect -1573 58 -1485 158
rect -1285 58 -497 158
rect -297 110 500 158
rect -297 58 697 110
rect 400 10 697 58
rect 897 10 994 110
<< polycont >>
rect 616 184 650 252
<< locali >>
rect -1806 512 -964 522
rect -1806 454 -1796 512
rect -1738 506 -964 512
rect -1738 466 -1730 506
rect -1040 466 -964 506
rect -1738 454 -964 466
rect -1806 450 -964 454
rect -1806 392 -1734 450
rect -1806 -176 -1790 392
rect -1750 -176 -1734 392
rect -1036 392 -964 450
rect 478 414 574 448
rect 1020 414 1116 448
rect -1036 252 -1020 392
rect -980 252 -964 392
rect -644 304 -620 338
rect -174 304 -150 338
rect 164 252 180 392
rect 220 252 236 392
rect 478 352 1116 414
rect 478 314 1082 352
rect 478 302 709 314
rect 693 280 709 302
rect 885 302 1082 314
rect 885 280 901 302
rect 616 252 650 268
rect -1477 209 -1461 243
rect -1309 209 -1293 243
rect -501 170 -485 204
rect -309 170 -293 204
rect 616 168 650 184
rect -501 12 -485 46
rect -309 12 -293 46
rect -1477 -27 -1461 7
rect -1309 -27 -1293 7
rect 693 -36 709 -2
rect 885 -36 901 -2
rect -1806 -234 -1734 -176
rect -1036 -176 -1020 -36
rect -980 -176 -964 -36
rect -644 -122 -620 -88
rect -174 -122 -150 -88
rect 164 -176 180 -36
rect 220 -176 236 -36
rect 1082 -136 1116 -74
rect 478 -170 574 -136
rect 1020 -170 1116 -136
rect -1036 -234 -964 -176
rect -1806 -250 -964 -234
rect -1806 -290 -1730 -250
rect -1040 -290 -964 -250
rect -1806 -306 -964 -290
<< viali >>
rect -1796 454 -1738 512
rect -1700 466 -1040 506
rect -1790 -176 -1750 392
rect 574 414 1020 448
rect -1020 252 -980 392
rect -620 304 -174 338
rect 180 252 220 392
rect 709 280 885 314
rect -1461 209 -1309 243
rect -485 170 -309 204
rect 616 184 650 252
rect 1082 194 1116 352
rect 1082 84 1116 194
rect -485 12 -309 46
rect -1461 -27 -1309 7
rect 709 -36 885 -2
rect -1020 -176 -980 -36
rect -620 -122 -174 -88
rect 180 -176 220 -36
rect 1082 -74 1116 84
rect 574 -170 1020 -136
rect -1730 -290 -1040 -250
<< metal1 >>
rect -1808 518 236 524
rect -1808 434 -1802 518
rect -1718 506 236 518
rect -1718 466 -1700 506
rect -1040 466 236 506
rect -1718 450 236 466
rect -1718 434 -1712 450
rect -1808 428 -1712 434
rect -1808 392 -1734 428
rect -1808 -176 -1790 392
rect -1750 -176 -1734 392
rect -1036 392 -964 450
rect -1036 252 -1020 392
rect -980 252 -964 392
rect 164 392 236 450
rect -632 338 -162 344
rect -632 304 -620 338
rect -174 304 -162 338
rect -632 298 -162 304
rect -1473 244 -1297 249
rect -1036 246 -964 252
rect -1473 243 -1454 244
rect -1316 243 -1297 244
rect -1473 209 -1461 243
rect -1309 209 -1297 243
rect -452 210 -352 298
rect 164 252 180 392
rect 220 252 236 392
rect 478 448 1122 454
rect 478 414 574 448
rect 1020 414 1122 448
rect 478 396 1122 414
rect 478 336 806 396
rect 696 314 806 336
rect 890 352 1122 396
rect 890 336 1082 352
rect 696 280 709 314
rect 890 312 898 336
rect 885 280 898 312
rect 696 274 898 280
rect -1473 203 -1454 209
rect -1461 192 -1454 203
rect -1316 203 -1297 209
rect -497 204 -297 210
rect -1316 192 -1309 203
rect -1461 24 -1309 192
rect -497 170 -485 204
rect -309 170 -297 204
rect -497 164 -297 170
rect -452 52 -352 164
rect -1461 13 -1454 24
rect -1473 7 -1454 13
rect -1316 13 -1309 24
rect -497 46 -297 52
rect -1316 7 -1297 13
rect -1473 -27 -1461 7
rect -1309 -27 -1297 7
rect -497 12 -485 46
rect -309 12 -297 46
rect -497 6 -297 12
rect -1473 -28 -1454 -27
rect -1316 -28 -1297 -27
rect -1473 -33 -1297 -28
rect -1808 -234 -1734 -176
rect -1036 -36 -964 -30
rect -1036 -176 -1020 -36
rect -980 -176 -964 -36
rect -452 -82 -352 6
rect 164 -36 236 252
rect 556 260 656 268
rect 556 176 564 260
rect 648 252 656 260
rect 650 184 656 252
rect 648 176 656 184
rect 556 168 656 176
rect -632 -88 -162 -82
rect -632 -122 -620 -88
rect -174 -122 -162 -88
rect -632 -128 -162 -122
rect -1036 -234 -964 -176
rect -1808 -250 -964 -234
rect -1808 -290 -1730 -250
rect -1040 -290 -964 -250
rect -1808 -306 -964 -290
rect -452 -204 -352 -128
rect 164 -176 180 -36
rect 220 -176 236 -36
rect 697 -2 897 4
rect 697 -36 709 -2
rect 885 -36 897 -2
rect 697 -42 756 -36
rect 748 -88 756 -42
rect 840 -42 897 -36
rect 840 -88 848 -42
rect 748 -96 848 -88
rect 1076 -74 1082 336
rect 1116 -74 1122 352
rect 1076 -130 1122 -74
rect 478 -136 1122 -130
rect 478 -170 574 -136
rect 1020 -170 1122 -136
rect 478 -176 1122 -170
rect 164 -182 236 -176
rect -452 -288 -444 -204
rect -360 -288 -352 -204
rect -452 -296 -352 -288
<< via1 >>
rect -1802 512 -1718 518
rect -1802 454 -1796 512
rect -1796 454 -1738 512
rect -1738 454 -1718 512
rect -1802 434 -1718 454
rect -1454 243 -1316 244
rect -1454 209 -1316 243
rect 806 314 890 396
rect 806 312 885 314
rect 885 312 890 314
rect -1454 192 -1316 209
rect -1454 7 -1316 24
rect -1454 -27 -1316 7
rect -1454 -28 -1316 -27
rect 564 252 648 260
rect 564 184 616 252
rect 616 184 648 252
rect 564 176 648 184
rect 756 -36 840 -4
rect 756 -88 840 -36
rect -444 -288 -360 -204
<< metal2 >>
rect -1810 518 -1710 526
rect -1810 434 -1802 518
rect -1718 434 -1710 518
rect -1810 426 -1710 434
rect 798 396 898 404
rect 798 312 806 396
rect 890 312 898 396
rect 798 304 898 312
rect 556 260 656 268
rect -1460 192 -1454 244
rect -1316 192 -1310 244
rect -1460 24 -1310 192
rect 556 176 564 260
rect 648 176 656 260
rect 556 168 656 176
rect -1460 -28 -1454 24
rect -1316 -28 -1310 24
rect 748 -4 848 4
rect 748 -88 756 -4
rect 840 -88 848 -4
rect 748 -96 848 -88
rect -452 -204 -352 -196
rect -452 -288 -444 -204
rect -360 -288 -352 -204
rect -452 -296 -352 -288
<< labels >>
flabel metal2 556 168 656 268 0 FreeSans 160 0 0 0 vinj_en_b
port 2 nsew signal input
flabel metal2 798 304 898 404 0 FreeSans 160 0 0 0 vinj
port 1 nsew power default
flabel metal2 748 -96 848 4 0 FreeSans 160 0 0 0 vsrc
port 5 nsew signal input
flabel metal2 -452 -296 -352 -196 0 FreeSans 160 0 0 0 vctrl
port 4 nsew analog input
flabel metal2 -1460 -28 -1310 244 0 FreeSans 160 0 0 0 vtun
port 3 nsew analog input
flabel metal2 -1810 426 -1710 526 0 FreeSans 160 0 0 0 VGND
port 6 nsew ground default
flabel poly -1154 58 -1054 158 0 FreeSans 160 0 0 0 fg
<< properties >>
string FIXED_BBOX -2010 -510 1394 726
<< end >>
