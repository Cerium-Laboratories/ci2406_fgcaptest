magic
tech sky130A
magscale 1 2
timestamp 1717562480
<< pwell >>
rect -284 -1582 284 1582
<< psubdiff >>
rect -248 1512 -152 1546
rect 152 1512 248 1546
rect -248 1450 -214 1512
rect 214 1450 248 1512
rect -248 -1512 -214 -1450
rect 214 -1512 248 -1450
rect -248 -1546 -152 -1512
rect 152 -1546 248 -1512
<< psubdiffcont >>
rect -152 1512 152 1546
rect -248 -1450 -214 1450
rect 214 -1450 248 1450
rect -152 -1546 152 -1512
<< xpolycontact >>
rect -118 984 -48 1416
rect -118 -1416 -48 -984
rect 48 984 118 1416
rect 48 -1416 118 -984
<< xpolyres >>
rect -118 -984 -48 984
rect 48 -984 118 984
<< locali >>
rect -248 1512 -152 1546
rect 152 1512 248 1546
rect -248 1450 -214 1512
rect 214 1450 248 1512
rect -248 -1512 -214 -1450
rect 214 -1512 248 -1450
rect -248 -1546 -152 -1512
rect 152 -1546 248 -1512
<< viali >>
rect -102 1001 -64 1398
rect 64 1001 102 1398
rect -102 -1398 -64 -1001
rect 64 -1398 102 -1001
<< metal1 >>
rect -108 1398 -58 1410
rect -108 1001 -102 1398
rect -64 1001 -58 1398
rect -108 989 -58 1001
rect 58 1398 108 1410
rect 58 1001 64 1398
rect 102 1001 108 1398
rect 58 989 108 1001
rect -108 -1001 -58 -989
rect -108 -1398 -102 -1001
rect -64 -1398 -58 -1001
rect -108 -1410 -58 -1398
rect 58 -1001 108 -989
rect 58 -1398 64 -1001
rect 102 -1398 108 -1001
rect 58 -1410 108 -1398
<< properties >>
string FIXED_BBOX -231 -1529 231 1529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
