magic
tech sky130A
magscale 1 2
timestamp 1717628967
<< poly >>
rect 2907 -5477 3240 -5380
rect 3140 -6470 3240 -5477
<< locali >>
rect 3076 -5154 3316 -5042
rect 3076 -5190 3282 -5154
<< metal1 >>
rect 3076 -5154 3322 -5036
rect 3276 -5190 3322 -5154
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3360 -5194 3460 -5188
rect 3502 -6650 3602 -6458
rect 3160 -6750 3602 -6650
rect 3140 -6812 3240 -6770
rect 3140 -6900 3146 -6812
rect 3234 -6900 3240 -6812
rect 3140 -6906 3240 -6900
rect 4006 -7030 4106 -5098
rect 2900 -7130 4106 -7030
<< via1 >>
rect 3366 -5188 3454 -5100
rect 3146 -6900 3234 -6812
<< metal2 >>
rect 3360 -5100 3460 -5094
rect 3360 -5188 3366 -5100
rect 3454 -5188 3460 -5100
rect 3360 -5222 3460 -5188
rect 2948 -5322 3460 -5222
rect 1294 -6812 3240 -6806
rect 1294 -6900 3146 -6812
rect 3234 -6900 3240 -6812
rect 1294 -6906 3240 -6900
use tg5v0  tg5v0_0
timestamp 1717628967
transform 0 -1 4094 1 0 -6628
box 28 0 1634 890
use fgcell  x1
timestamp 1717628967
transform 1 0 2010 0 1 -5490
box -1870 -310 1194 526
use diffamp_nmos  x2
timestamp 1717628967
transform 0 -1 3100 -1 0 -6070
box 20 -140 1140 2900
<< end >>
