magic
tech sky130A
timestamp 1717628967
<< psubdiff >>
rect 300 7228 6240 7240
rect 300 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 7116 6152 7128
rect 388 424 400 7116
rect 6140 424 6152 7116
rect 388 412 6152 424
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6240 7228
rect 300 300 6240 312
<< psubdiffcont >>
rect 312 312 388 7228
rect 440 7128 6100 7228
rect 440 312 6100 412
rect 6152 312 6228 7228
<< locali >>
rect 304 7228 6236 7236
rect 304 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 7120 6152 7128
rect 388 420 396 7120
rect 6144 420 6152 7120
rect 388 412 6152 420
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6236 7228
rect 304 304 6236 312
<< viali >>
rect 312 312 388 7228
rect 440 7128 6100 7228
rect 440 312 6100 412
rect 6152 312 6228 7228
<< metal1 >>
rect 304 7228 6236 7236
rect 304 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 7120 6152 7128
rect 388 420 396 7120
rect 6144 420 6152 7120
rect 388 412 6152 420
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6236 7228
rect 304 304 6236 312
<< via1 >>
rect 312 312 388 7228
rect 440 7128 6100 7228
rect 440 312 6100 412
rect 6152 312 6228 7228
<< metal2 >>
rect 304 7228 6236 7236
rect 304 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 7120 6152 7128
rect 388 420 396 7120
rect 6144 420 6152 7120
rect 388 412 6152 420
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6236 7228
rect 304 304 6236 312
<< via2 >>
rect 312 312 388 7228
rect 440 7128 6100 7228
rect 440 312 6100 412
rect 6152 312 6228 7228
<< metal3 >>
rect 304 7228 6236 7236
rect 304 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 7120 6152 7128
rect 388 420 396 7120
rect 6144 420 6152 7120
rect 388 412 6152 420
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6236 7228
rect 304 304 6236 312
<< via3 >>
rect 312 312 388 7228
rect 440 7128 6100 7228
rect 440 312 6100 412
rect 6152 312 6228 7228
<< metal4 >>
rect 270 7228 6270 7270
rect 270 312 312 7228
rect 388 7128 440 7228
rect 6100 7128 6152 7228
rect 388 412 6152 7128
rect 388 312 440 412
rect 6100 312 6152 412
rect 6228 312 6270 7228
rect 270 270 6270 312
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1717628967
transform 1 0 270 0 1 270
box -270 -270 6270 7270
<< end >>
