magic
tech sky130A
magscale 1 2
timestamp 1717034768
<< viali >>
rect 1132 -1053 1210 -975
rect 1132 -2621 1210 -2543
<< metal1 >>
rect 1126 -969 1216 -963
rect 1120 -1059 1126 -969
rect 1216 -1059 1222 -969
rect 1126 -1065 1216 -1059
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via1 >>
rect 1126 -975 1216 -969
rect 1126 -1053 1132 -975
rect 1132 -1053 1210 -975
rect 1210 -1053 1216 -975
rect 1126 -1059 1216 -1053
rect 1126 -2543 1216 -2537
rect 1126 -2621 1132 -2543
rect 1132 -2621 1210 -2543
rect 1210 -2621 1216 -2543
rect 1126 -2627 1216 -2621
<< metal2 >>
rect 1126 -969 1216 -963
rect 1122 -1054 1126 -974
rect 1216 -1054 1220 -974
rect 1126 -1065 1216 -1059
rect 1116 -2537 1226 -2532
rect 1116 -2627 1126 -2537
rect 1216 -2627 1226 -2537
rect 1116 -2632 1226 -2627
<< via2 >>
rect 1131 -1054 1211 -974
rect 1131 -2622 1211 -2542
<< metal3 >>
rect 1126 -974 1216 -963
rect 1126 -1054 1131 -974
rect 1211 -1054 1216 -974
rect 1126 -1682 1216 -1054
rect 1086 -1684 1356 -1682
rect 152 -1942 2208 -1684
rect 1126 -2538 1216 -2532
rect 1121 -2626 1127 -2538
rect 1215 -2626 1221 -2538
rect 1126 -2632 1216 -2626
<< via3 >>
rect 1127 -2542 1215 -2538
rect 1127 -2622 1131 -2542
rect 1131 -2622 1211 -2542
rect 1211 -2622 1215 -2542
rect 1127 -2626 1215 -2622
<< mimcap >>
rect 180 -1822 2180 -1712
rect 180 -1892 1136 -1822
rect 1206 -1892 2180 -1822
rect 180 -1914 2180 -1892
<< mimcapcontact >>
rect 1136 -1892 1206 -1822
<< metal4 >>
rect 1126 -1822 1216 -1812
rect 1126 -1892 1136 -1822
rect 1206 -1892 1216 -1822
rect 1126 -2538 1216 -1892
rect 1126 -2626 1127 -2538
rect 1215 -2626 1216 -2538
rect 1126 -2632 1216 -2626
use fgcell_amp  fgcell_amp_0 ~/Desktop/OpenCircuitDesign/ci2406_fgcaptest/mag
timestamp 1717034485
transform 1 0 -2 0 -1 -6399
box 2 -5898 6134 -3599
use fgcell_amp  fgcell_amp_1
timestamp 1717034485
transform 1 0 0 0 1 2800
box 2 -5898 6134 -3599
<< end >>
