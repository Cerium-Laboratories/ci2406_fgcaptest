magic
tech sky130A
magscale 1 2
timestamp 1717597427
<< error_s >>
rect 2764 -1602 3004 -1578
rect 2764 -1662 2788 -1602
rect 2980 -1662 3004 -1602
rect 2764 -1818 3004 -1662
rect 2460 -2038 2780 -1982
rect 884 -2282 1124 -2258
rect 884 -2474 908 -2282
rect 1100 -2474 1124 -2282
rect 2460 -2278 2484 -2038
rect 2700 -2278 2780 -2038
rect 4126 -2035 4214 -2030
rect 4126 -2113 4131 -2035
rect 4209 -2113 4214 -2035
rect 4126 -2118 4214 -2113
rect 2460 -2302 2780 -2278
rect 884 -2498 1124 -2474
rect 3334 -2487 3470 -2482
rect 3334 -2561 3339 -2487
rect 3465 -2561 3470 -2487
rect 3334 -2566 3470 -2561
rect 2862 -2625 3042 -2624
rect 2862 -2803 2863 -2625
rect 3041 -2803 3042 -2625
rect 2862 -2804 3042 -2803
rect 924 -3199 1104 -3198
rect 924 -3377 925 -3199
rect 1103 -3377 1104 -3199
rect 4258 -3202 4264 -3196
rect 4304 -3202 4310 -3196
rect 4252 -3208 4258 -3202
rect 4310 -3208 4316 -3202
rect 4252 -3254 4258 -3248
rect 4310 -3254 4316 -3248
rect 4258 -3260 4264 -3254
rect 4304 -3260 4310 -3254
rect 924 -3378 1104 -3377
rect 3786 -3390 3792 -3384
rect 3832 -3390 3838 -3384
rect 3780 -3396 3786 -3390
rect 3838 -3396 3844 -3390
rect 3780 -3442 3786 -3436
rect 3838 -3442 3844 -3436
rect 3786 -3448 3792 -3442
rect 3832 -3448 3838 -3442
rect 2764 -3902 3004 -3878
rect 2764 -4094 2788 -3902
rect 2980 -4094 3004 -3902
rect 2764 -4118 3004 -4094
<< polycont >>
rect 1526 -2400 1588 -2338
<< locali >>
rect 1510 -2331 1604 -2322
rect 1510 -2409 1516 -2331
rect 1594 -2409 1604 -2331
rect 1510 -2416 1604 -2409
<< viali >>
rect 1516 -2338 1594 -2331
rect 1516 -2400 1526 -2338
rect 1526 -2400 1588 -2338
rect 1588 -2400 1594 -2338
rect 1516 -2409 1594 -2400
<< metal1 >>
rect 2478 -2038 2730 -2028
rect 2478 -2278 2484 -2038
rect 2724 -2278 2730 -2038
rect 2478 -2284 2730 -2278
rect 1500 -2325 1610 -2320
rect 1500 -2415 1510 -2325
rect 1600 -2415 1610 -2325
rect 1500 -2420 1610 -2415
rect 4258 -3202 4316 -3196
rect 4310 -3254 4316 -3202
rect 4258 -3260 4316 -3254
rect 3780 -3390 3838 -3384
rect 3780 -3442 3786 -3390
rect 3780 -3448 3838 -3442
rect 786 -4020 1308 -4014
rect 1302 -4096 1308 -4020
rect 786 -4102 1308 -4096
<< via1 >>
rect 1660 -2020 1730 -1960
rect 2484 -2278 2724 -2038
rect 2884 -2178 3024 -2038
rect 4126 -2118 4214 -2030
rect 1510 -2331 1600 -2325
rect 1510 -2409 1516 -2331
rect 1516 -2409 1594 -2331
rect 1594 -2409 1600 -2331
rect 1510 -2415 1600 -2409
rect 4258 -3254 4310 -3202
rect 3786 -3442 3838 -3390
rect 786 -4096 1302 -4020
rect 2764 -4112 2944 -4024
<< metal2 >>
rect 1650 -1960 1740 -1954
rect 1650 -2020 1659 -1960
rect 1730 -2020 1740 -1960
rect 1650 -2028 1740 -2020
rect 2484 -2032 2724 -2028
rect 2478 -2038 2730 -2032
rect 878 -2258 1130 -2248
rect 878 -2498 884 -2258
rect 1124 -2498 1130 -2258
rect 2478 -2278 2484 -2038
rect 2724 -2278 2730 -2038
rect 2874 -2038 3034 -2028
rect 2874 -2178 2884 -2038
rect 3024 -2178 3034 -2038
rect 4116 -2030 4224 -2020
rect 4116 -2118 4126 -2030
rect 4214 -2118 4224 -2030
rect 4116 -2128 4224 -2118
rect 2874 -2188 3034 -2178
rect 2478 -2284 2730 -2278
rect 2484 -2288 2724 -2284
rect 1500 -2325 1610 -2320
rect 1500 -2415 1510 -2325
rect 1600 -2415 1610 -2325
rect 1500 -2420 1610 -2415
rect 878 -2508 1130 -2498
rect 3142 -2482 3480 -2472
rect 3142 -2566 3334 -2482
rect 3470 -2566 3480 -2482
rect 3142 -2576 3480 -2566
rect 914 -3912 1114 -3902
rect 914 -4014 924 -3912
rect 780 -4020 924 -4014
rect 1104 -4014 1114 -3912
rect 1104 -4020 1308 -4014
rect 780 -4096 786 -4020
rect 1302 -4096 1308 -4020
rect 780 -4102 1308 -4096
rect 2754 -4024 2954 -4018
rect 2754 -4112 2764 -4024
rect 2944 -4112 2954 -4024
rect 2754 -4118 2954 -4112
<< via2 >>
rect 1659 -2020 1660 -1960
rect 1660 -2020 1730 -1960
rect 884 -2498 1124 -2258
rect 2484 -2278 2724 -2038
rect 2884 -2178 3024 -2038
rect 4126 -2118 4214 -2030
rect 1515 -2410 1595 -2330
rect 3334 -2566 3470 -2482
rect 924 -4020 1104 -3912
rect 924 -4092 1104 -4020
rect 2764 -4112 2944 -4024
<< metal3 >>
rect 640 -1572 2720 -1560
rect 640 -1578 3010 -1572
rect 640 -1818 2764 -1578
rect 3004 -1818 3010 -1578
rect 640 -1824 3010 -1818
rect 640 -1840 2720 -1824
rect 1650 -1960 1740 -1840
rect 1650 -2020 1659 -1960
rect 1730 -2020 1740 -1960
rect 1650 -2030 1740 -2020
rect 2478 -2038 2730 -2032
rect 878 -2258 1130 -2252
rect 878 -2498 884 -2258
rect 1124 -2498 1130 -2258
rect 2478 -2278 2484 -2038
rect 2724 -2278 2730 -2038
rect 2478 -2284 2730 -2278
rect 2856 -2038 3048 -2028
rect 2856 -2178 2884 -2038
rect 3024 -2178 3048 -2038
rect 1510 -2326 1600 -2320
rect 1505 -2414 1511 -2326
rect 1599 -2414 1605 -2326
rect 1510 -2420 1600 -2414
rect 878 -2504 1130 -2498
rect 2856 -2624 3048 -2178
rect 2856 -2804 2862 -2624
rect 3042 -2804 3048 -2624
rect 2856 -2810 3048 -2804
rect 918 -3198 1110 -3192
rect 918 -3378 924 -3198
rect 1104 -3378 1110 -3198
rect 918 -3912 1110 -3378
rect 918 -4092 924 -3912
rect 1104 -4092 1110 -3912
rect 918 -4098 1110 -4092
rect 2758 -3938 2950 -3932
rect 2758 -4118 2764 -3938
rect 2944 -4118 2950 -3938
rect 2758 -4124 2950 -4118
<< via3 >>
rect 2764 -1818 3004 -1578
rect 884 -2498 1124 -2258
rect 2484 -2278 2724 -2038
rect 1511 -2330 1599 -2326
rect 1511 -2410 1515 -2330
rect 1515 -2410 1595 -2330
rect 1595 -2410 1599 -2330
rect 1511 -2414 1599 -2410
rect 2862 -2804 3042 -2624
rect 924 -3378 1104 -3198
rect 2764 -4024 2944 -3938
rect 2764 -4112 2944 -4024
rect 2764 -4118 2944 -4112
<< mimcap >>
rect 680 -1710 2680 -1600
rect 680 -1780 1520 -1710
rect 1590 -1780 2680 -1710
rect 680 -1800 2680 -1780
<< mimcapcontact >>
rect 1520 -1780 1590 -1710
<< metal4 >>
rect 2758 -1578 3010 -1572
rect 1510 -1710 1600 -1700
rect 1510 -1780 1520 -1710
rect 1590 -1780 1600 -1710
rect 878 -2258 1130 -2252
rect 878 -2498 884 -2258
rect 1124 -2498 1130 -2258
rect 1510 -2326 1600 -1780
rect 2758 -1818 2764 -1578
rect 3004 -1818 3010 -1578
rect 2758 -1824 3010 -1818
rect 2478 -2038 2730 -2032
rect 2478 -2278 2484 -2038
rect 2724 -2278 2730 -2038
rect 2478 -2284 2730 -2278
rect 1510 -2414 1511 -2326
rect 1599 -2414 1600 -2326
rect 1510 -2420 1600 -2414
rect 878 -2504 1130 -2498
rect 2758 -3878 3010 -3872
rect 2758 -4118 2764 -3878
rect 3004 -4118 3010 -3878
rect 2758 -4124 3010 -4118
<< via4 >>
rect 884 -2498 1124 -2258
rect 2764 -1818 3004 -1578
rect 2484 -2278 2724 -2038
rect 2764 -3938 3004 -3878
rect 2764 -4118 2944 -3938
rect 2944 -4118 3004 -3938
<< metal5 >>
rect 2460 -2038 2724 -1982
rect 2460 -2278 2484 -2038
rect 2460 -2302 2724 -2278
use fgcell_amp  x1
timestamp 1717597427
transform 1 0 384 0 1 3012
box 74 -7210 4106 -4964
<< labels >>
flabel via1 3786 -3442 3838 -3390 0 FreeSans 160 0 0 0 row_en
flabel via1 4258 -3254 4310 -3202 0 FreeSans 160 0 0 0 row_en_b
flabel via2 3334 -2566 3470 -2482 0 FreeSans 320 0 0 0 vsrc
flabel via3 2862 -2804 3042 -2624 0 FreeSans 320 0 0 0 vinj
flabel via3 924 -3378 1104 -3198 0 FreeSans 320 0 0 0 vdd
flabel via4 2764 -1818 3004 -1578 0 FreeSans 320 0 0 0 VGND
flabel via4 2484 -2278 2724 -2038 0 FreeSans 320 0 0 0 VGND
flabel via4 2764 -4118 3004 -3878 0 FreeSans 320 0 0 0 VGND
flabel via4 884 -2498 1124 -2258 0 FreeSans 480 0 0 0 vtun
<< end >>
