magic
tech sky130A
timestamp 1717628967
<< nwell >>
rect 1000 12515 1452 12605
rect 1000 11715 1452 11805
rect 1000 10915 1452 11005
rect 1000 10115 1452 10205
rect 1000 9315 1452 9405
rect 1000 8515 1452 8605
rect 1000 7715 1452 7805
rect 1000 6915 1452 7005
<< pwell >>
rect -1840 13220 -1790 13275
<< viali >>
rect -1765 13815 -1748 13852
rect -1766 13769 -1706 13786
rect -1765 13677 -1748 13737
rect -1766 13631 -1706 13648
rect -1765 13539 -1748 13599
rect -1766 13493 -1706 13510
rect -1765 13401 -1748 13461
rect -1766 13355 -1706 13372
rect -1098 13036 -1081 13053
rect -1028 13036 -1011 13053
rect -938 13000 -918 13080
rect -868 13036 -851 13053
rect -798 13036 -781 13053
rect -708 13000 -688 13080
rect -638 13036 -621 13053
rect -568 13036 -551 13053
rect -478 13000 -458 13080
rect -408 13036 -391 13053
rect -338 13036 -321 13053
rect -248 13000 -228 13080
rect -40 13036 -23 13053
rect 30 13036 47 13053
rect 120 13000 140 13080
rect 190 13036 207 13053
rect 260 13036 277 13053
rect 350 13000 370 13080
rect 420 13036 437 13053
rect 490 13036 507 13053
rect 580 13000 600 13080
rect 650 13036 667 13053
rect 720 13036 737 13053
rect 810 13000 830 13080
rect 1217 12806 1234 12823
rect 1355 12769 1372 12786
rect 1307 12731 1324 12748
rect 1355 12666 1372 12734
rect 1307 12372 1324 12389
rect 1355 12386 1372 12454
rect 1355 12334 1372 12351
rect 1217 12297 1234 12314
rect 1217 12006 1234 12023
rect 1355 11969 1372 11986
rect 1307 11931 1324 11948
rect 1355 11866 1372 11934
rect 1307 11572 1324 11589
rect 1355 11586 1372 11654
rect 1355 11534 1372 11551
rect 1217 11497 1234 11514
rect 1217 11206 1234 11223
rect 1355 11169 1372 11186
rect 1307 11131 1324 11148
rect 1355 11066 1372 11134
rect 1307 10772 1324 10789
rect 1355 10786 1372 10854
rect 1355 10734 1372 10751
rect 1217 10697 1234 10714
rect 1217 10406 1234 10423
rect 1355 10369 1372 10386
rect 1307 10331 1324 10348
rect 1355 10266 1372 10334
rect 1307 9972 1324 9989
rect 1355 9986 1372 10054
rect 1355 9934 1372 9951
rect 1217 9897 1234 9914
rect 1217 9606 1234 9623
rect 1355 9569 1372 9586
rect 1307 9531 1324 9548
rect 1355 9466 1372 9534
rect 1307 9172 1324 9189
rect 1355 9186 1372 9254
rect 1355 9134 1372 9151
rect 1217 9097 1234 9114
rect 1217 8806 1234 8823
rect 1355 8769 1372 8786
rect 1307 8731 1324 8748
rect 1355 8666 1372 8734
rect 1307 8372 1324 8389
rect 1355 8386 1372 8454
rect 1355 8334 1372 8351
rect 1217 8297 1234 8314
rect 1217 8006 1234 8023
rect 1355 7969 1372 7986
rect 1307 7931 1324 7948
rect 1355 7866 1372 7934
rect 1307 7572 1324 7589
rect 1355 7586 1372 7654
rect 1355 7534 1372 7551
rect 1217 7497 1234 7514
rect 1217 7206 1234 7223
rect 1355 7169 1372 7186
rect 1307 7131 1324 7148
rect 1355 7066 1372 7134
rect 1307 6772 1324 6789
rect 1355 6786 1372 6854
rect 1355 6734 1372 6751
rect 1217 6697 1234 6714
<< metal1 >>
rect -1772 13852 -1740 13857
rect -1772 13815 -1769 13852
rect -1743 13815 -1740 13852
rect -1564 13855 -817 13858
rect -1564 13829 -1561 13855
rect -1501 13829 -1102 13855
rect -1050 13829 -872 13855
rect -820 13829 -817 13855
rect -1564 13826 -817 13829
rect -1772 13809 -1740 13815
rect -1772 13786 -1700 13789
rect -1772 13760 -1766 13786
rect -1706 13760 -1700 13786
rect -1772 13757 -1700 13760
rect -1564 13786 -357 13789
rect -1564 13760 -1561 13786
rect -1501 13760 -642 13786
rect -590 13760 -412 13786
rect -360 13760 -357 13786
rect -1564 13757 -357 13760
rect -1772 13737 -1740 13743
rect -1772 13677 -1769 13737
rect -1743 13677 -1740 13737
rect -1564 13717 -517 13720
rect -1564 13691 -1561 13717
rect -1501 13691 -1032 13717
rect -980 13691 -572 13717
rect -520 13691 -517 13717
rect -1564 13688 -517 13691
rect -1772 13671 -1740 13677
rect -1772 13648 -1700 13651
rect -1772 13622 -1766 13648
rect -1706 13622 -1700 13648
rect -1772 13619 -1700 13622
rect -1564 13648 -287 13651
rect -1564 13622 -1561 13648
rect -1501 13622 -802 13648
rect -750 13622 -342 13648
rect -290 13622 -287 13648
rect -1564 13619 -287 13622
rect -1772 13599 -1740 13605
rect -1772 13539 -1769 13599
rect -1743 13539 -1740 13599
rect -1564 13579 241 13582
rect -1564 13553 -1561 13579
rect -1501 13553 -44 13579
rect 8 13553 186 13579
rect 238 13553 241 13579
rect -1564 13550 241 13553
rect -1772 13533 -1740 13539
rect -1772 13510 -1700 13513
rect -1772 13484 -1766 13510
rect -1706 13484 -1700 13510
rect -1772 13481 -1700 13484
rect -1564 13510 702 13513
rect -1564 13484 -1561 13510
rect -1501 13484 416 13510
rect 468 13484 646 13510
rect 698 13484 702 13510
rect -1564 13481 702 13484
rect -1772 13461 -1740 13467
rect -1772 13401 -1769 13461
rect -1743 13401 -1740 13461
rect -1564 13441 541 13444
rect -1564 13415 -1561 13441
rect -1501 13415 26 13441
rect 78 13415 486 13441
rect 538 13415 541 13441
rect -1564 13412 541 13415
rect -1772 13395 -1740 13401
rect -1772 13372 -1700 13375
rect -1772 13346 -1766 13372
rect -1706 13346 -1700 13372
rect -1772 13343 -1700 13346
rect -1564 13372 771 13375
rect -1564 13346 -1561 13372
rect -1501 13346 256 13372
rect 308 13346 716 13372
rect 768 13346 771 13372
rect -1564 13343 771 13346
rect -1900 12948 -1852 13273
rect -1628 13220 -1580 13273
rect -1628 13172 -1181 13220
rect 889 13217 1540 13220
rect 889 13172 933 13217
rect 930 13123 933 13172
rect 1427 13123 1540 13217
rect 930 13120 1540 13123
rect -941 13080 -915 13086
rect -1105 13031 -1102 13057
rect -1076 13031 -1073 13057
rect -1035 13031 -1032 13057
rect -1006 13031 -1003 13057
rect -711 13080 -685 13086
rect -875 13031 -872 13057
rect -846 13031 -843 13057
rect -805 13031 -802 13057
rect -776 13031 -773 13057
rect -941 12994 -915 13000
rect -481 13080 -455 13086
rect -645 13031 -642 13057
rect -616 13031 -613 13057
rect -575 13031 -572 13057
rect -546 13031 -543 13057
rect -711 12994 -685 13000
rect -251 13080 -225 13086
rect -415 13031 -412 13057
rect -386 13031 -383 13057
rect -345 13031 -342 13057
rect -316 13031 -313 13057
rect -481 12994 -455 13000
rect 117 13080 143 13086
rect -47 13031 -44 13057
rect -18 13031 -15 13057
rect 23 13031 26 13057
rect 52 13031 55 13057
rect -251 12994 -225 13000
rect 347 13080 373 13086
rect 183 13031 186 13057
rect 212 13031 215 13057
rect 253 13031 256 13057
rect 282 13031 285 13057
rect 117 12994 143 13000
rect 577 13080 603 13086
rect 413 13031 416 13057
rect 442 13031 445 13057
rect 483 13031 486 13057
rect 512 13031 515 13057
rect 347 12994 373 13000
rect 807 13080 833 13086
rect 643 13031 646 13057
rect 672 13031 675 13057
rect 713 13031 716 13057
rect 742 13031 745 13057
rect 577 12994 603 13000
rect 807 12994 833 13000
rect 930 13047 1433 13050
rect 930 12953 933 13047
rect 1427 12953 1433 13047
rect 930 12948 1433 12953
rect -1900 12945 -1181 12948
rect -1900 12904 -1237 12945
rect -1203 12904 -1181 12945
rect -1900 12900 -1181 12904
rect 889 12920 1433 12948
rect 889 12899 1019 12920
rect 798 12805 801 12831
rect 839 12826 842 12831
rect 839 12823 1240 12826
rect 839 12806 1217 12823
rect 1234 12806 1240 12823
rect 839 12805 1240 12806
rect 800 12803 1240 12805
rect -1242 12766 -1239 12792
rect -1201 12789 -1198 12792
rect -1201 12786 1378 12789
rect -1201 12769 1355 12786
rect 1372 12769 1378 12786
rect -1201 12766 1378 12769
rect -260 12725 -257 12751
rect -219 12748 1330 12751
rect -219 12731 1307 12748
rect 1324 12731 1330 12748
rect -219 12728 1330 12731
rect 1346 12734 1384 12737
rect -219 12725 -216 12728
rect 1346 12666 1352 12734
rect 1378 12666 1384 12734
rect 1346 12663 1384 12666
rect 1460 12600 1540 13120
rect 1019 12520 1540 12600
rect 1346 12454 1384 12457
rect -260 12369 -257 12395
rect -219 12392 -216 12395
rect -219 12389 1330 12392
rect -219 12372 1307 12389
rect 1324 12372 1330 12389
rect 1346 12386 1352 12454
rect 1378 12386 1384 12454
rect 1346 12383 1384 12386
rect -219 12369 1330 12372
rect -1242 12331 -1239 12357
rect -1201 12354 -1198 12357
rect -1201 12351 1378 12354
rect -1201 12334 1355 12351
rect 1372 12334 1378 12351
rect -1201 12331 1378 12334
rect 568 12291 571 12317
rect 609 12314 1240 12317
rect 609 12297 1217 12314
rect 1234 12297 1240 12314
rect 609 12294 1240 12297
rect 609 12291 612 12294
rect 930 12197 1433 12200
rect 930 12123 933 12197
rect 1007 12123 1433 12197
rect 930 12120 1433 12123
rect 338 12003 341 12029
rect 379 12026 382 12029
rect 379 12023 1240 12026
rect 379 12006 1217 12023
rect 1234 12006 1240 12023
rect 379 12003 1240 12006
rect -1242 11966 -1239 11992
rect -1201 11989 -1198 11992
rect -1201 11986 1378 11989
rect -1201 11969 1355 11986
rect 1372 11969 1378 11986
rect -1201 11966 1378 11969
rect -260 11925 -257 11951
rect -219 11948 1330 11951
rect -219 11931 1307 11948
rect 1324 11931 1330 11948
rect -219 11928 1330 11931
rect 1346 11934 1384 11937
rect -219 11925 -216 11928
rect 1346 11866 1352 11934
rect 1378 11866 1384 11934
rect 1346 11863 1384 11866
rect 1460 11800 1540 12520
rect 1019 11720 1540 11800
rect 1346 11654 1384 11657
rect -260 11572 -257 11598
rect -219 11592 -216 11598
rect -219 11589 1330 11592
rect -219 11572 1307 11589
rect 1324 11572 1330 11589
rect 1346 11586 1352 11654
rect 1378 11586 1384 11654
rect 1346 11583 1384 11586
rect -260 11569 1330 11572
rect -1242 11531 -1239 11557
rect -1201 11554 -1198 11557
rect -718 11554 -672 11560
rect -1201 11551 1378 11554
rect -1201 11534 1355 11551
rect 1372 11534 1378 11551
rect -1201 11531 1378 11534
rect 108 11491 111 11517
rect 149 11514 1240 11517
rect 149 11497 1217 11514
rect 1234 11497 1240 11514
rect 149 11494 1240 11497
rect 149 11491 152 11494
rect 930 11397 1433 11400
rect 930 11323 933 11397
rect 1007 11323 1433 11397
rect 930 11320 1433 11323
rect 798 11205 801 11231
rect 839 11226 842 11231
rect 839 11223 1240 11226
rect 839 11206 1217 11223
rect 1234 11206 1240 11223
rect 839 11205 1240 11206
rect 800 11203 1240 11205
rect -1242 11166 -1239 11192
rect -1201 11189 -1198 11192
rect -1201 11186 1378 11189
rect -1201 11169 1355 11186
rect 1372 11169 1378 11186
rect -1201 11166 1378 11169
rect -490 11125 -487 11151
rect -449 11148 1330 11151
rect -449 11131 1307 11148
rect 1324 11131 1330 11148
rect -449 11128 1330 11131
rect 1346 11134 1384 11137
rect -449 11125 -446 11128
rect 1346 11066 1352 11134
rect 1378 11066 1384 11134
rect 1346 11063 1384 11066
rect 1460 11000 1540 11720
rect 1019 10920 1540 11000
rect 1346 10854 1384 10857
rect -490 10769 -487 10795
rect -449 10792 -446 10795
rect -449 10789 1330 10792
rect -449 10772 1307 10789
rect 1324 10772 1330 10789
rect 1346 10786 1352 10854
rect 1378 10786 1384 10854
rect 1346 10783 1384 10786
rect -449 10769 1330 10772
rect -1242 10731 -1239 10757
rect -1201 10754 -1198 10757
rect -1201 10751 1378 10754
rect -1201 10734 1355 10751
rect 1372 10734 1378 10751
rect -1201 10731 1378 10734
rect 568 10691 571 10717
rect 609 10714 1240 10717
rect 609 10697 1217 10714
rect 1234 10697 1240 10714
rect 609 10694 1240 10697
rect 609 10691 612 10694
rect 930 10597 1433 10600
rect 930 10523 933 10597
rect 1007 10523 1433 10597
rect 930 10520 1433 10523
rect 338 10403 341 10429
rect 379 10426 382 10429
rect 379 10423 1240 10426
rect 379 10406 1217 10423
rect 1234 10406 1240 10423
rect 379 10403 1240 10406
rect -1242 10366 -1239 10392
rect -1201 10389 -1198 10392
rect -1201 10386 1378 10389
rect -1201 10369 1355 10386
rect 1372 10369 1378 10386
rect -1201 10366 1378 10369
rect -490 10325 -487 10351
rect -449 10348 1330 10351
rect -449 10331 1307 10348
rect 1324 10331 1330 10348
rect -449 10328 1330 10331
rect 1346 10334 1384 10337
rect -449 10325 -446 10328
rect 1346 10266 1352 10334
rect 1378 10266 1384 10334
rect 1346 10263 1384 10266
rect 1460 10200 1540 10920
rect 1019 10120 1540 10200
rect 1346 10054 1384 10057
rect -490 9998 -446 9999
rect -490 9972 -487 9998
rect -449 9992 -446 9998
rect -449 9989 1330 9992
rect -449 9972 1307 9989
rect 1324 9972 1330 9989
rect 1346 9986 1352 10054
rect 1378 9986 1384 10054
rect 1346 9983 1384 9986
rect -490 9969 1330 9972
rect -490 9968 -446 9969
rect -1242 9931 -1239 9957
rect -1201 9954 -1198 9957
rect -1201 9951 1378 9954
rect -1201 9934 1355 9951
rect 1372 9934 1378 9951
rect -1201 9931 1378 9934
rect 108 9891 111 9917
rect 149 9914 1240 9917
rect 149 9897 1217 9914
rect 1234 9897 1240 9914
rect 149 9894 1240 9897
rect 149 9891 152 9894
rect 930 9797 1433 9800
rect 930 9723 933 9797
rect 1007 9723 1433 9797
rect 930 9720 1433 9723
rect 798 9605 801 9631
rect 839 9626 842 9631
rect 839 9623 1240 9626
rect 839 9606 1217 9623
rect 1234 9606 1240 9623
rect 839 9605 1240 9606
rect 800 9603 1240 9605
rect -1242 9566 -1239 9592
rect -1201 9589 -1198 9592
rect -1201 9586 1378 9589
rect -1201 9569 1355 9586
rect 1372 9569 1378 9586
rect -1201 9566 1378 9569
rect -717 9525 -714 9551
rect -676 9548 1330 9551
rect -676 9531 1307 9548
rect 1324 9531 1330 9548
rect -676 9528 1330 9531
rect 1346 9534 1384 9537
rect -676 9525 -673 9528
rect 1346 9466 1352 9534
rect 1378 9466 1384 9534
rect 1346 9463 1384 9466
rect 1460 9400 1540 10120
rect 1019 9320 1540 9400
rect 1346 9254 1384 9257
rect -717 9169 -714 9195
rect -676 9192 -673 9195
rect -676 9189 1330 9192
rect -676 9172 1307 9189
rect 1324 9172 1330 9189
rect 1346 9186 1352 9254
rect 1378 9186 1384 9254
rect 1346 9183 1384 9186
rect -676 9169 1330 9172
rect -1242 9131 -1239 9157
rect -1201 9154 -1198 9157
rect -1201 9151 1378 9154
rect -1201 9134 1355 9151
rect 1372 9134 1378 9151
rect -1201 9131 1378 9134
rect 568 9091 571 9117
rect 609 9114 1240 9117
rect 609 9097 1217 9114
rect 1234 9097 1240 9114
rect 609 9094 1240 9097
rect 609 9091 612 9094
rect 930 8997 1433 9000
rect 930 8923 933 8997
rect 1007 8923 1433 8997
rect 930 8920 1433 8923
rect 338 8803 341 8829
rect 379 8826 382 8829
rect 379 8823 1240 8826
rect 379 8806 1217 8823
rect 1234 8806 1240 8823
rect 379 8803 1240 8806
rect -1242 8766 -1239 8792
rect -1201 8789 -1198 8792
rect -1201 8786 1378 8789
rect -1201 8769 1355 8786
rect 1372 8769 1378 8786
rect -1201 8766 1378 8769
rect -717 8725 -714 8751
rect -676 8748 1330 8751
rect -676 8731 1307 8748
rect 1324 8731 1330 8748
rect -676 8728 1330 8731
rect 1346 8734 1384 8737
rect -676 8725 -673 8728
rect 1346 8666 1352 8734
rect 1378 8666 1384 8734
rect 1346 8663 1384 8666
rect 1460 8600 1540 9320
rect 1019 8520 1540 8600
rect 1346 8454 1384 8457
rect -717 8398 -673 8399
rect -717 8371 -714 8398
rect -676 8392 -673 8398
rect -676 8389 1330 8392
rect -676 8372 1307 8389
rect 1324 8372 1330 8389
rect 1346 8386 1352 8454
rect 1378 8386 1384 8454
rect 1346 8383 1384 8386
rect -676 8371 1330 8372
rect -717 8369 1330 8371
rect -1242 8331 -1239 8357
rect -1201 8354 -1198 8357
rect -1201 8351 1378 8354
rect -1201 8334 1355 8351
rect 1372 8334 1378 8351
rect -1201 8331 1378 8334
rect 108 8291 111 8317
rect 149 8314 1240 8317
rect 149 8297 1217 8314
rect 1234 8297 1240 8314
rect 149 8294 1240 8297
rect 149 8291 152 8294
rect 930 8197 1433 8200
rect 930 8123 933 8197
rect 1007 8123 1433 8197
rect 930 8120 1433 8123
rect 798 8005 801 8031
rect 839 8026 842 8031
rect 839 8023 1240 8026
rect 839 8006 1217 8023
rect 1234 8006 1240 8023
rect 839 8005 1240 8006
rect 798 8003 1240 8005
rect -1242 7966 -1239 7992
rect -1201 7989 -1198 7992
rect -1201 7986 1378 7989
rect -1201 7969 1355 7986
rect 1372 7969 1378 7986
rect -1201 7966 1378 7969
rect -950 7925 -947 7951
rect -909 7948 1330 7951
rect -909 7931 1307 7948
rect 1324 7931 1330 7948
rect -909 7928 1330 7931
rect 1346 7934 1384 7937
rect -909 7925 -906 7928
rect 1346 7866 1352 7934
rect 1378 7866 1384 7934
rect 1346 7863 1384 7866
rect 1460 7800 1540 8520
rect 1019 7720 1540 7800
rect 1346 7654 1384 7657
rect -950 7569 -947 7595
rect -909 7592 -906 7595
rect -909 7589 1330 7592
rect -909 7572 1307 7589
rect 1324 7572 1330 7589
rect 1346 7586 1352 7654
rect 1378 7586 1384 7654
rect 1346 7583 1384 7586
rect -909 7569 1330 7572
rect -1242 7531 -1239 7557
rect -1201 7554 -1198 7557
rect -1201 7551 1378 7554
rect -1201 7534 1355 7551
rect 1372 7534 1378 7551
rect -1201 7531 1378 7534
rect 568 7491 571 7517
rect 609 7514 1240 7517
rect 609 7497 1217 7514
rect 1234 7497 1240 7514
rect 609 7494 1240 7497
rect 609 7491 612 7494
rect 930 7397 1433 7400
rect 930 7323 933 7397
rect 1007 7323 1433 7397
rect 930 7320 1433 7323
rect 338 7203 341 7229
rect 379 7226 382 7229
rect 379 7223 1240 7226
rect 379 7206 1217 7223
rect 1234 7206 1240 7223
rect 379 7203 1240 7206
rect -1242 7166 -1239 7192
rect -1201 7189 -1198 7192
rect -1201 7186 1378 7189
rect -1201 7169 1355 7186
rect 1372 7169 1378 7186
rect -1201 7166 1378 7169
rect -950 7125 -947 7151
rect -909 7148 1330 7151
rect -909 7131 1307 7148
rect 1324 7131 1330 7148
rect -909 7128 1330 7131
rect 1346 7134 1384 7137
rect -909 7125 -906 7128
rect 1346 7066 1352 7134
rect 1378 7066 1384 7134
rect 1346 7063 1384 7066
rect 1460 7000 1540 7720
rect 1019 6920 1540 7000
rect 1346 6854 1384 6857
rect -950 6800 -906 6803
rect -950 6774 -948 6800
rect -908 6792 -906 6800
rect -908 6789 1330 6792
rect -908 6774 1307 6789
rect -950 6772 1307 6774
rect 1324 6772 1330 6789
rect 1346 6786 1352 6854
rect 1378 6786 1384 6854
rect 1346 6783 1384 6786
rect -950 6769 1330 6772
rect -1242 6731 -1239 6757
rect -1201 6754 -1198 6757
rect -1201 6751 1378 6754
rect -1201 6734 1355 6751
rect 1372 6734 1378 6751
rect -1201 6731 1378 6734
rect -1242 6728 -1198 6731
rect 108 6691 111 6717
rect 149 6714 1240 6717
rect 149 6697 1217 6714
rect 1234 6697 1240 6714
rect 149 6694 1240 6697
rect 149 6691 152 6694
rect 108 6688 152 6691
rect 930 6597 1433 6600
rect 930 6523 933 6597
rect 1007 6523 1433 6597
rect 930 6520 1433 6523
<< via1 >>
rect -1769 13815 -1765 13852
rect -1765 13815 -1748 13852
rect -1748 13815 -1743 13852
rect -1561 13829 -1501 13855
rect -1102 13829 -1050 13855
rect -872 13829 -820 13855
rect -1766 13769 -1706 13786
rect -1766 13760 -1706 13769
rect -1561 13760 -1501 13786
rect -642 13760 -590 13786
rect -412 13760 -360 13786
rect -1769 13677 -1765 13737
rect -1765 13677 -1748 13737
rect -1748 13677 -1743 13737
rect -1561 13691 -1501 13717
rect -1032 13691 -980 13717
rect -572 13691 -520 13717
rect -1766 13631 -1706 13648
rect -1766 13622 -1706 13631
rect -1561 13622 -1501 13648
rect -802 13622 -750 13648
rect -342 13622 -290 13648
rect -1769 13539 -1765 13599
rect -1765 13539 -1748 13599
rect -1748 13539 -1743 13599
rect -1561 13553 -1501 13579
rect -44 13553 8 13579
rect 186 13553 238 13579
rect -1766 13493 -1706 13510
rect -1766 13484 -1706 13493
rect -1561 13484 -1501 13510
rect 416 13484 468 13510
rect 646 13484 698 13510
rect -1769 13401 -1765 13461
rect -1765 13401 -1748 13461
rect -1748 13401 -1743 13461
rect -1561 13415 -1501 13441
rect 26 13415 78 13441
rect 486 13415 538 13441
rect -1766 13355 -1706 13372
rect -1766 13346 -1706 13355
rect -1561 13346 -1501 13372
rect 256 13346 308 13372
rect 716 13346 768 13372
rect 933 13123 1427 13217
rect -1102 13053 -1076 13057
rect -1102 13036 -1098 13053
rect -1098 13036 -1081 13053
rect -1081 13036 -1076 13053
rect -1102 13031 -1076 13036
rect -1032 13053 -1006 13057
rect -1032 13036 -1028 13053
rect -1028 13036 -1011 13053
rect -1011 13036 -1006 13053
rect -1032 13031 -1006 13036
rect -941 13000 -938 13080
rect -938 13000 -918 13080
rect -918 13000 -915 13080
rect -872 13053 -846 13057
rect -872 13036 -868 13053
rect -868 13036 -851 13053
rect -851 13036 -846 13053
rect -872 13031 -846 13036
rect -802 13053 -776 13057
rect -802 13036 -798 13053
rect -798 13036 -781 13053
rect -781 13036 -776 13053
rect -802 13031 -776 13036
rect -711 13000 -708 13080
rect -708 13000 -688 13080
rect -688 13000 -685 13080
rect -642 13053 -616 13057
rect -642 13036 -638 13053
rect -638 13036 -621 13053
rect -621 13036 -616 13053
rect -642 13031 -616 13036
rect -572 13053 -546 13057
rect -572 13036 -568 13053
rect -568 13036 -551 13053
rect -551 13036 -546 13053
rect -572 13031 -546 13036
rect -481 13000 -478 13080
rect -478 13000 -458 13080
rect -458 13000 -455 13080
rect -412 13053 -386 13057
rect -412 13036 -408 13053
rect -408 13036 -391 13053
rect -391 13036 -386 13053
rect -412 13031 -386 13036
rect -342 13053 -316 13057
rect -342 13036 -338 13053
rect -338 13036 -321 13053
rect -321 13036 -316 13053
rect -342 13031 -316 13036
rect -251 13000 -248 13080
rect -248 13000 -228 13080
rect -228 13000 -225 13080
rect -44 13053 -18 13057
rect -44 13036 -40 13053
rect -40 13036 -23 13053
rect -23 13036 -18 13053
rect -44 13031 -18 13036
rect 26 13053 52 13057
rect 26 13036 30 13053
rect 30 13036 47 13053
rect 47 13036 52 13053
rect 26 13031 52 13036
rect 117 13000 120 13080
rect 120 13000 140 13080
rect 140 13000 143 13080
rect 186 13053 212 13057
rect 186 13036 190 13053
rect 190 13036 207 13053
rect 207 13036 212 13053
rect 186 13031 212 13036
rect 256 13053 282 13057
rect 256 13036 260 13053
rect 260 13036 277 13053
rect 277 13036 282 13053
rect 256 13031 282 13036
rect 347 13000 350 13080
rect 350 13000 370 13080
rect 370 13000 373 13080
rect 416 13053 442 13057
rect 416 13036 420 13053
rect 420 13036 437 13053
rect 437 13036 442 13053
rect 416 13031 442 13036
rect 486 13053 512 13057
rect 486 13036 490 13053
rect 490 13036 507 13053
rect 507 13036 512 13053
rect 486 13031 512 13036
rect 577 13000 580 13080
rect 580 13000 600 13080
rect 600 13000 603 13080
rect 646 13053 672 13057
rect 646 13036 650 13053
rect 650 13036 667 13053
rect 667 13036 672 13053
rect 646 13031 672 13036
rect 716 13053 742 13057
rect 716 13036 720 13053
rect 720 13036 737 13053
rect 737 13036 742 13053
rect 716 13031 742 13036
rect 807 13000 810 13080
rect 810 13000 830 13080
rect 830 13000 833 13080
rect 933 12953 1427 13047
rect -1237 12904 -1203 12945
rect 801 12805 839 12831
rect -1239 12766 -1201 12792
rect -257 12725 -219 12751
rect 1352 12666 1355 12734
rect 1355 12666 1372 12734
rect 1372 12666 1378 12734
rect -257 12369 -219 12395
rect 1352 12386 1355 12454
rect 1355 12386 1372 12454
rect 1372 12386 1378 12454
rect -1239 12331 -1201 12357
rect 571 12291 609 12317
rect 933 12123 1007 12197
rect 341 12003 379 12029
rect -1239 11966 -1201 11992
rect -257 11925 -219 11951
rect 1352 11866 1355 11934
rect 1355 11866 1372 11934
rect 1372 11866 1378 11934
rect -257 11572 -219 11598
rect 1352 11586 1355 11654
rect 1355 11586 1372 11654
rect 1372 11586 1378 11654
rect -1239 11531 -1201 11557
rect 111 11491 149 11517
rect 933 11323 1007 11397
rect 801 11205 839 11231
rect -1239 11166 -1201 11192
rect -487 11125 -449 11151
rect 1352 11066 1355 11134
rect 1355 11066 1372 11134
rect 1372 11066 1378 11134
rect -487 10769 -449 10795
rect 1352 10786 1355 10854
rect 1355 10786 1372 10854
rect 1372 10786 1378 10854
rect -1239 10731 -1201 10757
rect 571 10691 609 10717
rect 933 10523 1007 10597
rect 341 10403 379 10429
rect -1239 10366 -1201 10392
rect -487 10325 -449 10351
rect 1352 10266 1355 10334
rect 1355 10266 1372 10334
rect 1372 10266 1378 10334
rect -487 9972 -449 9998
rect 1352 9986 1355 10054
rect 1355 9986 1372 10054
rect 1372 9986 1378 10054
rect -1239 9931 -1201 9957
rect 111 9891 149 9917
rect 933 9723 1007 9797
rect 801 9605 839 9631
rect -1239 9566 -1201 9592
rect -714 9525 -676 9551
rect 1352 9466 1355 9534
rect 1355 9466 1372 9534
rect 1372 9466 1378 9534
rect -714 9169 -676 9195
rect 1352 9186 1355 9254
rect 1355 9186 1372 9254
rect 1372 9186 1378 9254
rect -1239 9131 -1201 9157
rect 571 9091 609 9117
rect 933 8923 1007 8997
rect 341 8803 379 8829
rect -1239 8766 -1201 8792
rect -714 8725 -676 8751
rect 1352 8666 1355 8734
rect 1355 8666 1372 8734
rect 1372 8666 1378 8734
rect -714 8371 -676 8398
rect 1352 8386 1355 8454
rect 1355 8386 1372 8454
rect 1372 8386 1378 8454
rect -1239 8331 -1201 8357
rect 111 8291 149 8317
rect 933 8123 1007 8197
rect 801 8005 839 8031
rect -1239 7966 -1201 7992
rect -947 7925 -909 7951
rect 1352 7866 1355 7934
rect 1355 7866 1372 7934
rect 1372 7866 1378 7934
rect -947 7569 -909 7595
rect 1352 7586 1355 7654
rect 1355 7586 1372 7654
rect 1372 7586 1378 7654
rect -1239 7531 -1201 7557
rect 571 7491 609 7517
rect 933 7323 1007 7397
rect 341 7203 379 7229
rect -1239 7166 -1201 7192
rect -947 7125 -909 7151
rect 1352 7066 1355 7134
rect 1355 7066 1372 7134
rect 1372 7066 1378 7134
rect -948 6774 -908 6800
rect 1352 6786 1355 6854
rect 1355 6786 1372 6854
rect 1372 6786 1378 6854
rect -1239 6731 -1201 6757
rect 111 6691 149 6717
rect 933 6523 1007 6597
<< metal2 >>
rect -2020 13878 -1920 13902
rect -2020 13852 -1900 13878
rect -1580 13855 -1498 13858
rect -1580 13852 -1561 13855
rect -2020 13815 -1769 13852
rect -1743 13829 -1561 13852
rect -1501 13829 -1498 13855
rect -1743 13826 -1498 13829
rect -1105 13855 -1047 13858
rect -1105 13829 -1102 13855
rect -1050 13829 -1047 13855
rect -1105 13826 -1047 13829
rect -875 13855 -817 13858
rect -875 13829 -872 13855
rect -820 13829 -817 13855
rect -875 13826 -817 13829
rect -1743 13815 -1740 13826
rect -2020 13812 -1740 13815
rect -2020 13802 -1920 13812
rect -1769 13786 -1498 13789
rect -2020 13740 -1920 13764
rect -1769 13760 -1766 13786
rect -1706 13760 -1561 13786
rect -1501 13760 -1498 13786
rect -1769 13757 -1498 13760
rect -2020 13737 -1740 13740
rect -2020 13677 -1769 13737
rect -1743 13720 -1740 13737
rect -1743 13717 -1498 13720
rect -1743 13691 -1561 13717
rect -1501 13691 -1498 13717
rect -1743 13688 -1498 13691
rect -1743 13677 -1740 13688
rect -2020 13674 -1740 13677
rect -2020 13664 -1920 13674
rect -1769 13648 -1498 13651
rect -2020 13602 -1920 13626
rect -1769 13622 -1766 13648
rect -1706 13622 -1561 13648
rect -1501 13622 -1498 13648
rect -1769 13619 -1498 13622
rect -2020 13599 -1740 13602
rect -2020 13539 -1769 13599
rect -1743 13582 -1740 13599
rect -1743 13579 -1498 13582
rect -1743 13553 -1561 13579
rect -1501 13553 -1498 13579
rect -1743 13550 -1498 13553
rect -1743 13539 -1740 13550
rect -2020 13536 -1740 13539
rect -2020 13526 -1920 13536
rect -1769 13510 -1498 13513
rect -2020 13464 -1920 13488
rect -1769 13484 -1766 13510
rect -1706 13484 -1561 13510
rect -1501 13484 -1498 13510
rect -1769 13481 -1498 13484
rect -2020 13461 -1740 13464
rect -2020 13401 -1769 13461
rect -1743 13444 -1740 13461
rect -1743 13441 -1498 13444
rect -1743 13415 -1561 13441
rect -1501 13415 -1498 13441
rect -1743 13412 -1498 13415
rect -1743 13401 -1740 13412
rect -2020 13398 -1740 13401
rect -2020 13388 -1920 13398
rect -1769 13372 -1498 13375
rect -1769 13346 -1766 13372
rect -1706 13346 -1561 13372
rect -1501 13346 -1498 13372
rect -1769 13343 -1498 13346
rect -1105 13057 -1073 13826
rect -1105 13031 -1102 13057
rect -1076 13031 -1073 13057
rect -1105 13028 -1073 13031
rect -1035 13717 -977 13720
rect -1035 13691 -1032 13717
rect -980 13691 -977 13717
rect -1035 13688 -977 13691
rect -1035 13057 -1003 13688
rect -1035 13031 -1032 13057
rect -1006 13031 -1003 13057
rect -1035 13028 -1003 13031
rect -948 13080 -908 13090
rect -948 13000 -941 13080
rect -915 13000 -908 13080
rect -875 13057 -843 13826
rect -645 13786 -587 13789
rect -645 13760 -642 13786
rect -590 13760 -587 13786
rect -645 13757 -587 13760
rect -415 13786 -357 13789
rect -415 13760 -412 13786
rect -360 13760 -357 13786
rect -415 13757 -357 13760
rect -875 13031 -872 13057
rect -846 13031 -843 13057
rect -875 13028 -843 13031
rect -805 13648 -747 13651
rect -805 13622 -802 13648
rect -750 13622 -747 13648
rect -805 13619 -747 13622
rect -805 13057 -773 13619
rect -805 13031 -802 13057
rect -776 13031 -773 13057
rect -805 13028 -773 13031
rect -715 13080 -675 13094
rect -1240 12945 -1200 12948
rect -1240 12904 -1237 12945
rect -1203 12904 -1200 12945
rect -1240 12792 -1200 12904
rect -1240 12766 -1239 12792
rect -1201 12766 -1200 12792
rect -1240 12357 -1200 12766
rect -1240 12331 -1239 12357
rect -1201 12331 -1200 12357
rect -1240 11992 -1200 12331
rect -1240 11966 -1239 11992
rect -1201 11966 -1200 11992
rect -1240 11557 -1200 11966
rect -1240 11531 -1239 11557
rect -1201 11531 -1200 11557
rect -1240 11192 -1200 11531
rect -1240 11166 -1239 11192
rect -1201 11166 -1200 11192
rect -1240 10757 -1200 11166
rect -1240 10731 -1239 10757
rect -1201 10731 -1200 10757
rect -1240 10392 -1200 10731
rect -1240 10366 -1239 10392
rect -1201 10366 -1200 10392
rect -1240 9957 -1200 10366
rect -1240 9931 -1239 9957
rect -1201 9931 -1200 9957
rect -1240 9592 -1200 9931
rect -1240 9566 -1239 9592
rect -1201 9566 -1200 9592
rect -1240 9157 -1200 9566
rect -1240 9131 -1239 9157
rect -1201 9131 -1200 9157
rect -1240 8792 -1200 9131
rect -1240 8766 -1239 8792
rect -1201 8766 -1200 8792
rect -1240 8357 -1200 8766
rect -1240 8331 -1239 8357
rect -1201 8331 -1200 8357
rect -1240 7992 -1200 8331
rect -1240 7966 -1239 7992
rect -1201 7966 -1200 7992
rect -1240 7557 -1200 7966
rect -1240 7531 -1239 7557
rect -1201 7531 -1200 7557
rect -1240 7192 -1200 7531
rect -1240 7166 -1239 7192
rect -1201 7166 -1200 7192
rect -1240 6757 -1200 7166
rect -948 7951 -908 13000
rect -715 13000 -711 13080
rect -685 13000 -675 13080
rect -645 13057 -613 13757
rect -645 13031 -642 13057
rect -616 13031 -613 13057
rect -645 13028 -613 13031
rect -575 13717 -517 13720
rect -575 13691 -572 13717
rect -520 13691 -517 13717
rect -575 13688 -517 13691
rect -575 13057 -543 13688
rect -575 13031 -572 13057
rect -546 13031 -543 13057
rect -575 13028 -543 13031
rect -488 13080 -448 13090
rect -715 9551 -675 13000
rect -488 13000 -481 13080
rect -455 13000 -448 13080
rect -415 13057 -383 13757
rect -415 13031 -412 13057
rect -386 13031 -383 13057
rect -415 13028 -383 13031
rect -345 13648 -287 13651
rect -345 13622 -342 13648
rect -290 13622 -287 13648
rect -345 13619 -287 13622
rect -345 13057 -313 13619
rect -47 13579 11 13582
rect -47 13553 -44 13579
rect 8 13553 11 13579
rect -47 13550 11 13553
rect 183 13579 241 13582
rect 183 13553 186 13579
rect 238 13553 241 13579
rect 183 13550 241 13553
rect -345 13031 -342 13057
rect -316 13031 -313 13057
rect -345 13028 -313 13031
rect -258 13080 -218 13090
rect -488 11151 -448 13000
rect -258 13000 -251 13080
rect -225 13000 -218 13080
rect -47 13057 -15 13550
rect -47 13031 -44 13057
rect -18 13031 -15 13057
rect -47 13028 -15 13031
rect 23 13441 81 13444
rect 23 13415 26 13441
rect 78 13415 81 13441
rect 23 13412 81 13415
rect 23 13057 55 13412
rect 23 13031 26 13057
rect 52 13031 55 13057
rect 23 13028 55 13031
rect 110 13080 150 13090
rect -258 12751 -218 13000
rect -258 12725 -257 12751
rect -219 12725 -218 12751
rect -258 12395 -218 12725
rect -258 12369 -257 12395
rect -219 12369 -218 12395
rect -258 11951 -218 12369
rect -258 11925 -257 11951
rect -219 11925 -218 11951
rect -258 11598 -218 11925
rect 110 13000 117 13080
rect 143 13000 150 13080
rect 183 13057 215 13550
rect 413 13510 471 13513
rect 413 13484 416 13510
rect 468 13484 471 13510
rect 413 13481 471 13484
rect 643 13510 701 13513
rect 643 13484 646 13510
rect 698 13484 701 13510
rect 643 13481 701 13484
rect 183 13031 186 13057
rect 212 13031 215 13057
rect 183 13028 215 13031
rect 253 13372 311 13375
rect 253 13346 256 13372
rect 308 13346 311 13372
rect 253 13343 311 13346
rect 253 13057 285 13343
rect 253 13031 256 13057
rect 282 13031 285 13057
rect 253 13028 285 13031
rect 340 13080 380 13090
rect -260 11572 -257 11598
rect -219 11572 -216 11598
rect -260 11569 -216 11572
rect -488 11125 -487 11151
rect -449 11125 -448 11151
rect -488 10795 -448 11125
rect -488 10769 -487 10795
rect -449 10769 -448 10795
rect -488 10351 -448 10769
rect -488 10325 -487 10351
rect -449 10325 -448 10351
rect -488 9998 -448 10325
rect -488 9972 -487 9998
rect -449 9972 -448 9998
rect -488 9969 -448 9972
rect 110 11517 150 13000
rect 110 11491 111 11517
rect 149 11491 150 11517
rect -715 9525 -714 9551
rect -676 9525 -675 9551
rect -715 9195 -675 9525
rect -715 9169 -714 9195
rect -676 9169 -675 9195
rect -715 8751 -675 9169
rect -715 8725 -714 8751
rect -676 8725 -675 8751
rect -715 8399 -675 8725
rect 110 9917 150 11491
rect 110 9891 111 9917
rect 149 9891 150 9917
rect -717 8398 -673 8399
rect -717 8371 -714 8398
rect -676 8371 -673 8398
rect -717 8369 -673 8371
rect -948 7925 -947 7951
rect -909 7925 -908 7951
rect -948 7595 -908 7925
rect -948 7569 -947 7595
rect -909 7569 -908 7595
rect -948 7151 -908 7569
rect -948 7125 -947 7151
rect -909 7125 -908 7151
rect -948 6803 -908 7125
rect 110 8317 150 9891
rect 110 8291 111 8317
rect 149 8291 150 8317
rect -950 6800 -906 6803
rect -950 6774 -948 6800
rect -908 6774 -906 6800
rect -950 6769 -906 6774
rect -1242 6731 -1239 6757
rect -1201 6731 -1198 6757
rect -1242 6728 -1198 6731
rect 110 6718 150 8291
rect 340 13000 347 13080
rect 373 13000 380 13080
rect 413 13057 445 13481
rect 413 13031 416 13057
rect 442 13031 445 13057
rect 413 13028 445 13031
rect 483 13441 541 13444
rect 483 13415 486 13441
rect 538 13415 541 13441
rect 483 13412 541 13415
rect 483 13057 515 13412
rect 483 13031 486 13057
rect 512 13031 515 13057
rect 483 13028 515 13031
rect 570 13080 610 13090
rect 340 12029 380 13000
rect 340 12003 341 12029
rect 379 12003 380 12029
rect 340 10429 380 12003
rect 340 10403 341 10429
rect 379 10403 380 10429
rect 340 8829 380 10403
rect 340 8803 341 8829
rect 379 8803 380 8829
rect 340 7234 380 8803
rect 570 13000 577 13080
rect 603 13000 610 13080
rect 643 13057 675 13481
rect 643 13031 646 13057
rect 672 13031 675 13057
rect 643 13028 675 13031
rect 713 13372 771 13375
rect 713 13346 716 13372
rect 768 13346 771 13372
rect 713 13343 771 13346
rect 713 13057 745 13343
rect 930 13217 1430 13220
rect 930 13123 933 13217
rect 1427 13123 1430 13217
rect 930 13120 1430 13123
rect 713 13031 716 13057
rect 742 13031 745 13057
rect 713 13028 745 13031
rect 800 13080 840 13090
rect 570 12317 610 13000
rect 570 12291 571 12317
rect 609 12291 610 12317
rect 570 10717 610 12291
rect 570 10691 571 10717
rect 609 10691 610 10717
rect 570 9117 610 10691
rect 570 9091 571 9117
rect 609 9091 610 9117
rect 570 7517 610 9091
rect 800 13000 807 13080
rect 833 13000 840 13080
rect 800 12831 840 13000
rect 800 12805 801 12831
rect 839 12805 840 12831
rect 800 11231 840 12805
rect 800 11205 801 11231
rect 839 11205 840 11231
rect 800 9631 840 11205
rect 800 9605 801 9631
rect 839 9605 840 9631
rect 800 8031 840 9605
rect 930 13047 1430 13050
rect 930 12953 933 13047
rect 1427 12953 1430 13047
rect 930 12950 1430 12953
rect 930 12197 1010 12950
rect 1460 12737 1560 12800
rect 1349 12734 1560 12737
rect 1349 12666 1352 12734
rect 1378 12700 1560 12734
rect 1378 12666 1381 12700
rect 1349 12663 1381 12666
rect 1349 12454 1381 12457
rect 1349 12386 1352 12454
rect 1378 12400 1381 12454
rect 1378 12386 1560 12400
rect 1349 12363 1560 12386
rect 1460 12300 1560 12363
rect 930 12123 933 12197
rect 1007 12123 1010 12197
rect 930 11397 1010 12123
rect 1460 11937 1560 12000
rect 1349 11934 1560 11937
rect 1349 11866 1352 11934
rect 1378 11900 1560 11934
rect 1378 11866 1381 11900
rect 1349 11863 1381 11866
rect 1349 11654 1381 11657
rect 1349 11586 1352 11654
rect 1378 11600 1381 11654
rect 1378 11586 1560 11600
rect 1349 11563 1560 11586
rect 1460 11500 1560 11563
rect 930 11323 933 11397
rect 1007 11323 1010 11397
rect 930 10597 1010 11323
rect 1460 11137 1560 11200
rect 1349 11134 1560 11137
rect 1349 11066 1352 11134
rect 1378 11100 1560 11134
rect 1378 11066 1381 11100
rect 1349 11063 1381 11066
rect 1349 10854 1381 10857
rect 1349 10786 1352 10854
rect 1378 10800 1381 10854
rect 1378 10786 1560 10800
rect 1349 10763 1560 10786
rect 1460 10700 1560 10763
rect 930 10523 933 10597
rect 1007 10523 1010 10597
rect 930 9797 1010 10523
rect 1460 10337 1560 10400
rect 1349 10334 1560 10337
rect 1349 10266 1352 10334
rect 1378 10300 1560 10334
rect 1378 10266 1381 10300
rect 1349 10263 1381 10266
rect 1349 10054 1381 10057
rect 1349 9986 1352 10054
rect 1378 10000 1381 10054
rect 1378 9986 1560 10000
rect 1349 9963 1560 9986
rect 1460 9900 1560 9963
rect 930 9723 933 9797
rect 1007 9723 1010 9797
rect 930 8997 1010 9723
rect 1460 9537 1560 9600
rect 1349 9534 1560 9537
rect 1349 9466 1352 9534
rect 1378 9500 1560 9534
rect 1378 9466 1381 9500
rect 1349 9463 1381 9466
rect 1349 9254 1381 9257
rect 1349 9186 1352 9254
rect 1378 9200 1381 9254
rect 1378 9186 1560 9200
rect 1349 9163 1560 9186
rect 1460 9100 1560 9163
rect 930 8923 933 8997
rect 1007 8923 1010 8997
rect 930 8197 1010 8923
rect 1460 8737 1560 8800
rect 1349 8734 1560 8737
rect 1349 8666 1352 8734
rect 1378 8700 1560 8734
rect 1378 8666 1381 8700
rect 1349 8663 1381 8666
rect 1349 8454 1381 8457
rect 1349 8386 1352 8454
rect 1378 8400 1381 8454
rect 1378 8386 1560 8400
rect 1349 8363 1560 8386
rect 1460 8300 1560 8363
rect 930 8123 933 8197
rect 1007 8123 1010 8197
rect 798 8005 801 8031
rect 839 8005 842 8031
rect 798 8003 842 8005
rect 570 7491 571 7517
rect 609 7491 610 7517
rect 570 7488 610 7491
rect 338 7229 380 7234
rect 338 7203 341 7229
rect 379 7203 380 7229
rect 338 7200 380 7203
rect 930 7397 1010 8123
rect 1460 7937 1560 8000
rect 1349 7934 1560 7937
rect 1349 7866 1352 7934
rect 1378 7900 1560 7934
rect 1378 7866 1381 7900
rect 1349 7863 1381 7866
rect 1349 7654 1381 7657
rect 1349 7586 1352 7654
rect 1378 7600 1381 7654
rect 1378 7586 1560 7600
rect 1349 7563 1560 7586
rect 1460 7500 1560 7563
rect 930 7323 933 7397
rect 1007 7323 1010 7397
rect 108 6717 152 6718
rect 108 6691 111 6717
rect 149 6691 152 6717
rect 108 6689 152 6691
rect 930 6597 1010 7323
rect 1460 7137 1560 7200
rect 1349 7134 1560 7137
rect 1349 7066 1352 7134
rect 1378 7100 1560 7134
rect 1378 7066 1381 7100
rect 1349 7063 1381 7066
rect 1349 6854 1381 6857
rect 1349 6786 1352 6854
rect 1378 6800 1381 6854
rect 1378 6786 1560 6800
rect 1349 6763 1560 6786
rect 1460 6700 1560 6763
rect 930 6523 933 6597
rect 1007 6523 1010 6597
rect 930 6520 1010 6523
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
array 0 0 -452 0 7 -800
timestamp 1717628967
transform -1 0 1203 0 -1 7296
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
array 0 0 452 0 7 800
timestamp 1717628967
transform 1 0 1066 0 1 6624
box -19 -24 157 296
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1717628967
transform 1 0 -215 0 1 12924
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717628967
transform 1 0 383 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
array 0 0 -452 0 7 -800
timestamp 1717628967
transform -1 0 1387 0 -1 7296
box -19 -24 203 296
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_1
array 0 0 -452 0 7 800
timestamp 1717628967
transform -1 0 1388 0 1 6624
box -19 -24 203 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
array 0 0 -452 0 7 -800
timestamp 1717628967
transform -1 0 1433 0 -1 7296
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
array 0 0 -452 0 7 -800
timestamp 1717628967
transform -1 0 1065 0 -1 7296
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
array 0 0 452 0 7 800
timestamp 1717628967
transform 1 0 1020 0 1 6624
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
array 0 0 452 0 7 800
timestamp 1717628967
transform 1 0 1388 0 1 6624
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1717628967
transform 1 0 -1181 0 1 12924
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1717628967
transform 1 0 843 0 1 12924
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1717628967
transform 0 1 -1876 -1 0 13917
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1717628967
transform 0 1 -1876 -1 0 13319
box -19 -24 65 296
use sky130_fd_sc_hd__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717628967
transform 0 1 -1876 -1 0 13871
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x3
timestamp 1717628967
transform 0 1 -1876 -1 0 13733
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x4
timestamp 1717628967
transform 0 1 -1876 -1 0 13595
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x5
timestamp 1717628967
transform 0 1 -1876 -1 0 13457
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_2  x6
timestamp 1717628967
transform 1 0 613 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x8
timestamp 1717628967
transform 1 0 153 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x9
timestamp 1717628967
transform 1 0 -77 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x10
timestamp 1717628967
transform 1 0 -445 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x11
timestamp 1717628967
transform 1 0 -675 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x12
timestamp 1717628967
transform 1 0 -905 0 1 12924
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_2  x13
timestamp 1717628967
transform 1 0 -1135 0 1 12924
box -19 -24 249 296
<< labels >>
flabel metal2 1460 7100 1560 7200 0 FreeSans 160 0 0 0 w[14]
port 24 nsew
flabel metal2 1460 7500 1560 7600 0 FreeSans 160 0 0 0 w[13]
port 25 nsew
flabel metal2 1460 7900 1560 8000 0 FreeSans 160 0 0 0 w[12]
port 26 nsew
flabel metal2 1460 8300 1560 8400 0 FreeSans 160 0 0 0 w[11]
port 27 nsew
flabel metal2 1460 8700 1560 8800 0 FreeSans 160 0 0 0 w[10]
port 28 nsew
flabel metal2 1460 9100 1560 9200 0 FreeSans 160 0 0 0 w[9]
port 29 nsew
flabel metal2 1460 9500 1560 9600 0 FreeSans 160 0 0 0 w[8]
port 30 nsew
flabel metal2 1460 9900 1560 10000 0 FreeSans 160 0 0 0 w[7]
port 31 nsew
flabel metal2 1460 10300 1560 10400 0 FreeSans 160 0 0 0 w[6]
port 32 nsew
flabel metal2 1460 10700 1560 10800 0 FreeSans 160 0 0 0 w[5]
port 33 nsew
flabel metal2 1460 11100 1560 11200 0 FreeSans 160 0 0 0 w[4]
port 34 nsew
flabel metal2 1460 11500 1560 11600 0 FreeSans 160 0 0 0 w[3]
port 35 nsew
flabel metal2 1460 11900 1560 12000 0 FreeSans 160 0 0 0 w[2]
port 36 nsew
flabel metal2 1460 12300 1560 12400 0 FreeSans 160 0 0 0 w[1]
port 37 nsew
flabel metal2 -2020 13802 -1920 13902 0 FreeSans 160 0 0 0 a[3]
port 3 nsew
flabel metal2 -2020 13664 -1920 13764 0 FreeSans 160 0 0 0 a[2]
port 4 nsew
flabel metal2 -2020 13526 -1920 13626 0 FreeSans 160 0 0 0 a[1]
port 5 nsew
flabel metal2 -2020 13388 -1920 13488 0 FreeSans 160 0 0 0 a[0]
port 6 nsew
flabel metal2 1460 12700 1560 12800 0 FreeSans 160 0 0 0 w[0]
port 38 nsew
flabel metal2 1330 12950 1430 13050 0 FreeSans 160 0 0 0 VGND
port 1 nsew
flabel metal2 1330 13120 1430 13220 0 FreeSans 160 0 0 0 VPWR
port 0 nsew
flabel pwell -1840 13220 -1790 13270 0 FreeSans 160 0 0 0 VGND
flabel metal2 1460 6700 1560 6800 0 FreeSans 160 0 0 0 w[15]
port 23 nsew
<< end >>
