magic
tech sky130A
timestamp 1716945357
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vout
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 v1
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 v2
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 vb
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 VDD
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 VSS
port 5 nsew
<< end >>
